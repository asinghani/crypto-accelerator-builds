magic
tech sky130A
magscale 1 2
timestamp 1608101209
<< locali >>
rect 8125 685899 8159 695453
rect 72525 684607 72559 694093
rect 137845 685899 137879 695453
rect 219081 685899 219115 695453
rect 72801 676107 72835 684437
rect 154313 676243 154347 685797
rect 218989 666587 219023 676141
rect 72985 647275 73019 656829
rect 219265 647275 219299 656829
rect 73077 616879 73111 626501
rect 219357 616879 219391 626501
rect 219081 608719 219115 611405
rect 219265 601579 219299 608549
rect 72893 589339 72927 598893
rect 219173 589339 219207 598893
rect 8033 579751 8067 589237
rect 137753 579751 137787 589237
rect 154313 579751 154347 589237
rect 72617 569959 72651 579581
rect 137569 569959 137603 579581
rect 218897 569959 218931 579581
rect 72617 550647 72651 553401
rect 137661 550647 137695 560201
rect 218897 550647 218931 553401
rect 8033 540991 8067 550545
rect 72617 531335 72651 534089
rect 154405 521679 154439 531233
rect 154405 502367 154439 511921
rect 7941 444431 7975 453985
rect 154221 444431 154255 453985
rect 163513 162911 163547 172465
rect 188077 169303 188111 173961
rect 220093 173655 220127 173825
rect 221749 173043 221783 173757
rect 229385 172907 229419 173213
rect 229477 172567 229511 173553
rect 229569 172635 229603 173349
rect 229661 173247 229695 173485
rect 229753 173315 229787 173553
rect 299489 173315 299523 173485
rect 309057 173383 309091 173485
rect 229845 172771 229879 173281
rect 234537 173043 234571 173281
rect 239321 172907 239355 173145
rect 299489 173043 299523 173145
rect 304273 173043 304307 173145
rect 239413 172703 239447 172873
rect 354597 172839 354631 173213
rect 163053 151827 163087 161381
rect 181177 145027 181211 162809
rect 206017 154615 206051 164169
rect 223865 162911 223899 172465
rect 225337 151827 225371 161381
rect 240517 156315 240551 164169
rect 385233 157335 385267 164169
rect 157625 124219 157659 133841
rect 159005 131019 159039 143497
rect 163145 128299 163179 143497
rect 179613 134555 179647 143497
rect 181085 134011 181119 143497
rect 181085 124219 181119 133841
rect 183845 124287 183879 143497
rect 207305 128299 207339 143497
rect 210065 128299 210099 135201
rect 219633 134011 219667 143497
rect 223773 142171 223807 151725
rect 240425 133943 240459 138125
rect 385233 137955 385267 144857
rect 158913 113203 158947 122757
rect 158913 103547 158947 113033
rect 163145 108987 163179 115889
rect 181177 114563 181211 115957
rect 180993 104907 181027 114393
rect 183937 113203 183971 122757
rect 196173 115991 196207 125545
rect 197645 115991 197679 125545
rect 222393 124219 222427 133841
rect 223773 122859 223807 124253
rect 218345 114563 218379 119357
rect 219633 114563 219667 119357
rect 185133 111027 185167 114461
rect 228097 106335 228131 115889
rect 240425 114563 240459 124117
rect 385049 106335 385083 119357
rect 158913 85595 158947 95081
rect 163145 89675 163179 96577
rect 174185 95251 174219 104805
rect 182465 103615 182499 104873
rect 182557 97291 182591 102085
rect 196173 96679 196207 106233
rect 197645 96679 197679 106233
rect 218253 100011 218287 104737
rect 217057 96611 217091 99433
rect 181085 85595 181119 95149
rect 174185 75939 174219 85493
rect 183845 84235 183879 85765
rect 185041 85595 185075 95149
rect 218253 91851 218287 95149
rect 219541 92463 219575 98685
rect 222485 96679 222519 106233
rect 240425 96679 240459 106233
rect 385049 93891 385083 104805
rect 182465 79339 182499 84133
rect 209881 77299 209915 86921
rect 219449 82875 219483 92429
rect 228005 82875 228039 92429
rect 181085 66283 181119 75837
rect 183845 66283 183879 70669
rect 207121 70363 207155 77197
rect 219633 75939 219667 82841
rect 159005 56627 159039 66181
rect 180993 57919 181027 60809
rect 180993 46971 181027 56525
rect 182373 48331 182407 64821
rect 183845 55267 183879 64821
rect 185225 59211 185259 64821
rect 193505 48331 193539 57885
rect 210065 48331 210099 57885
rect 216965 56627 216999 67541
rect 222485 63563 222519 73117
rect 228005 64923 228039 77945
rect 239045 77299 239079 86921
rect 240425 77299 240459 86921
rect 256893 67643 256927 77197
rect 237297 56627 237331 66181
rect 238677 56627 238711 66181
rect 240425 62747 240459 67541
rect 385049 66283 385083 84133
rect 218253 46971 218287 56525
rect 158913 29087 158947 46869
rect 163145 29019 163179 38573
rect 182373 37315 182407 46869
rect 210065 37315 210099 46869
rect 181085 29019 181119 34697
rect 182373 29019 182407 31705
rect 156429 12427 156463 19261
rect 158913 19227 158947 27557
rect 181177 18003 181211 27557
rect 183753 26367 183787 27693
rect 207397 27659 207431 37213
rect 219541 35955 219575 38709
rect 221013 37315 221047 46869
rect 222577 45611 222611 54621
rect 239045 48331 239079 57885
rect 237297 37315 237331 46869
rect 238677 37315 238711 46869
rect 239045 37315 239079 38709
rect 385325 29019 385359 38573
rect 183753 16643 183787 26197
rect 183753 8075 183787 13141
rect 185133 4335 185167 12461
rect 200405 9707 200439 19261
rect 207213 18003 207247 22117
rect 216965 9707 216999 27557
rect 219541 9707 219575 27557
rect 226625 19975 226659 28917
rect 222485 11747 222519 19261
rect 237205 9707 237239 27489
rect 238401 9707 238435 27489
rect 239045 22763 239079 28917
rect 257077 12291 257111 19261
rect 385049 9707 385083 19261
rect 42809 3315 42843 3485
rect 84761 3179 84795 4029
rect 84853 3383 84887 4029
rect 93777 3179 93811 4097
rect 167009 3655 167043 3757
rect 162133 3451 162167 3621
rect 170597 3655 170631 3825
rect 162041 3383 162075 3417
rect 162225 3383 162259 3621
rect 174001 3587 174035 3689
rect 162041 3349 162259 3383
rect 111073 3213 111935 3247
rect 111073 3179 111107 3213
rect 107669 2839 107703 3145
rect 111809 3043 111843 3145
rect 111901 3043 111935 3213
rect 121503 2873 121653 2907
rect 107519 2805 107703 2839
rect 201417 1887 201451 3621
rect 202889 3519 202923 3621
rect 206109 1275 206143 3553
rect 211169 3519 211203 3757
rect 220093 3723 220127 3961
rect 220737 3519 220771 3757
rect 222209 3043 222243 5797
rect 224877 3451 224911 3757
rect 226441 3587 226475 3893
rect 229511 3825 229753 3859
rect 226349 3043 226383 3553
rect 230489 3519 230523 4777
rect 234721 3995 234755 4097
rect 234629 3723 234663 3961
rect 304825 3689 306297 3723
rect 304825 3655 304859 3689
rect 233525 3043 233559 3485
rect 243001 3247 243035 3417
rect 275661 3383 275695 3621
rect 306147 3553 306297 3587
rect 319913 2975 319947 3145
rect 320005 3009 320557 3043
rect 320005 2907 320039 3009
rect 325433 2907 325467 3077
rect 255053 595 255087 2805
<< viali >>
rect 8125 695453 8159 695487
rect 137845 695453 137879 695487
rect 8125 685865 8159 685899
rect 72525 694093 72559 694127
rect 137845 685865 137879 685899
rect 219081 695453 219115 695487
rect 219081 685865 219115 685899
rect 72525 684573 72559 684607
rect 154313 685797 154347 685831
rect 72801 684437 72835 684471
rect 154313 676209 154347 676243
rect 72801 676073 72835 676107
rect 218989 676141 219023 676175
rect 218989 666553 219023 666587
rect 72985 656829 73019 656863
rect 72985 647241 73019 647275
rect 219265 656829 219299 656863
rect 219265 647241 219299 647275
rect 73077 626501 73111 626535
rect 73077 616845 73111 616879
rect 219357 626501 219391 626535
rect 219357 616845 219391 616879
rect 219081 611405 219115 611439
rect 219081 608685 219115 608719
rect 219265 608549 219299 608583
rect 219265 601545 219299 601579
rect 72893 598893 72927 598927
rect 72893 589305 72927 589339
rect 219173 598893 219207 598927
rect 219173 589305 219207 589339
rect 8033 589237 8067 589271
rect 8033 579717 8067 579751
rect 137753 589237 137787 589271
rect 137753 579717 137787 579751
rect 154313 589237 154347 589271
rect 154313 579717 154347 579751
rect 72617 579581 72651 579615
rect 72617 569925 72651 569959
rect 137569 579581 137603 579615
rect 137569 569925 137603 569959
rect 218897 579581 218931 579615
rect 218897 569925 218931 569959
rect 137661 560201 137695 560235
rect 72617 553401 72651 553435
rect 72617 550613 72651 550647
rect 137661 550613 137695 550647
rect 218897 553401 218931 553435
rect 218897 550613 218931 550647
rect 8033 550545 8067 550579
rect 8033 540957 8067 540991
rect 72617 534089 72651 534123
rect 72617 531301 72651 531335
rect 154405 531233 154439 531267
rect 154405 521645 154439 521679
rect 154405 511921 154439 511955
rect 154405 502333 154439 502367
rect 7941 453985 7975 454019
rect 7941 444397 7975 444431
rect 154221 453985 154255 454019
rect 154221 444397 154255 444431
rect 188077 173961 188111 173995
rect 163513 172465 163547 172499
rect 220093 173825 220127 173859
rect 220093 173621 220127 173655
rect 221749 173757 221783 173791
rect 229477 173553 229511 173587
rect 221749 173009 221783 173043
rect 229385 173213 229419 173247
rect 229385 172873 229419 172907
rect 229753 173553 229787 173587
rect 229661 173485 229695 173519
rect 229569 173349 229603 173383
rect 299489 173485 299523 173519
rect 309057 173485 309091 173519
rect 309057 173349 309091 173383
rect 229753 173281 229787 173315
rect 229845 173281 229879 173315
rect 229661 173213 229695 173247
rect 234537 173281 234571 173315
rect 299489 173281 299523 173315
rect 354597 173213 354631 173247
rect 234537 173009 234571 173043
rect 239321 173145 239355 173179
rect 299489 173145 299523 173179
rect 299489 173009 299523 173043
rect 304273 173145 304307 173179
rect 304273 173009 304307 173043
rect 239321 172873 239355 172907
rect 239413 172873 239447 172907
rect 229845 172737 229879 172771
rect 354597 172805 354631 172839
rect 239413 172669 239447 172703
rect 229569 172601 229603 172635
rect 229477 172533 229511 172567
rect 188077 169269 188111 169303
rect 223865 172465 223899 172499
rect 163513 162877 163547 162911
rect 206017 164169 206051 164203
rect 181177 162809 181211 162843
rect 163053 161381 163087 161415
rect 163053 151793 163087 151827
rect 223865 162877 223899 162911
rect 240517 164169 240551 164203
rect 206017 154581 206051 154615
rect 225337 161381 225371 161415
rect 385233 164169 385267 164203
rect 385233 157301 385267 157335
rect 240517 156281 240551 156315
rect 225337 151793 225371 151827
rect 181177 144993 181211 145027
rect 223773 151725 223807 151759
rect 159005 143497 159039 143531
rect 157625 133841 157659 133875
rect 159005 130985 159039 131019
rect 163145 143497 163179 143531
rect 179613 143497 179647 143531
rect 179613 134521 179647 134555
rect 181085 143497 181119 143531
rect 181085 133977 181119 134011
rect 183845 143497 183879 143531
rect 163145 128265 163179 128299
rect 181085 133841 181119 133875
rect 157625 124185 157659 124219
rect 207305 143497 207339 143531
rect 219633 143497 219667 143531
rect 207305 128265 207339 128299
rect 210065 135201 210099 135235
rect 223773 142137 223807 142171
rect 385233 144857 385267 144891
rect 219633 133977 219667 134011
rect 240425 138125 240459 138159
rect 385233 137921 385267 137955
rect 240425 133909 240459 133943
rect 210065 128265 210099 128299
rect 222393 133841 222427 133875
rect 183845 124253 183879 124287
rect 196173 125545 196207 125579
rect 181085 124185 181119 124219
rect 158913 122757 158947 122791
rect 183937 122757 183971 122791
rect 181177 115957 181211 115991
rect 158913 113169 158947 113203
rect 163145 115889 163179 115923
rect 158913 113033 158947 113067
rect 181177 114529 181211 114563
rect 163145 108953 163179 108987
rect 180993 114393 181027 114427
rect 196173 115957 196207 115991
rect 197645 125545 197679 125579
rect 222393 124185 222427 124219
rect 223773 124253 223807 124287
rect 223773 122825 223807 122859
rect 240425 124117 240459 124151
rect 197645 115957 197679 115991
rect 218345 119357 218379 119391
rect 218345 114529 218379 114563
rect 219633 119357 219667 119391
rect 219633 114529 219667 114563
rect 228097 115889 228131 115923
rect 183937 113169 183971 113203
rect 185133 114461 185167 114495
rect 185133 110993 185167 111027
rect 240425 114529 240459 114563
rect 385049 119357 385083 119391
rect 228097 106301 228131 106335
rect 385049 106301 385083 106335
rect 196173 106233 196207 106267
rect 180993 104873 181027 104907
rect 182465 104873 182499 104907
rect 158913 103513 158947 103547
rect 174185 104805 174219 104839
rect 163145 96577 163179 96611
rect 158913 95081 158947 95115
rect 182465 103581 182499 103615
rect 182557 102085 182591 102119
rect 182557 97257 182591 97291
rect 196173 96645 196207 96679
rect 197645 106233 197679 106267
rect 222485 106233 222519 106267
rect 218253 104737 218287 104771
rect 218253 99977 218287 100011
rect 197645 96645 197679 96679
rect 217057 99433 217091 99467
rect 217057 96577 217091 96611
rect 219541 98685 219575 98719
rect 174185 95217 174219 95251
rect 163145 89641 163179 89675
rect 181085 95149 181119 95183
rect 158913 85561 158947 85595
rect 185041 95149 185075 95183
rect 181085 85561 181119 85595
rect 183845 85765 183879 85799
rect 174185 85493 174219 85527
rect 218253 95149 218287 95183
rect 222485 96645 222519 96679
rect 240425 106233 240459 106267
rect 240425 96645 240459 96679
rect 385049 104805 385083 104839
rect 385049 93857 385083 93891
rect 218253 91817 218287 91851
rect 219449 92429 219483 92463
rect 219541 92429 219575 92463
rect 228005 92429 228039 92463
rect 185041 85561 185075 85595
rect 209881 86921 209915 86955
rect 183845 84201 183879 84235
rect 182465 84133 182499 84167
rect 182465 79305 182499 79339
rect 219449 82841 219483 82875
rect 219633 82841 219667 82875
rect 228005 82841 228039 82875
rect 239045 86921 239079 86955
rect 209881 77265 209915 77299
rect 174185 75905 174219 75939
rect 207121 77197 207155 77231
rect 181085 75837 181119 75871
rect 181085 66249 181119 66283
rect 183845 70669 183879 70703
rect 219633 75905 219667 75939
rect 228005 77945 228039 77979
rect 207121 70329 207155 70363
rect 222485 73117 222519 73151
rect 183845 66249 183879 66283
rect 216965 67541 216999 67575
rect 159005 66181 159039 66215
rect 182373 64821 182407 64855
rect 180993 60809 181027 60843
rect 180993 57885 181027 57919
rect 159005 56593 159039 56627
rect 180993 56525 181027 56559
rect 183845 64821 183879 64855
rect 185225 64821 185259 64855
rect 185225 59177 185259 59211
rect 183845 55233 183879 55267
rect 193505 57885 193539 57919
rect 182373 48297 182407 48331
rect 193505 48297 193539 48331
rect 210065 57885 210099 57919
rect 239045 77265 239079 77299
rect 240425 86921 240459 86955
rect 240425 77265 240459 77299
rect 385049 84133 385083 84167
rect 256893 77197 256927 77231
rect 256893 67609 256927 67643
rect 240425 67541 240459 67575
rect 228005 64889 228039 64923
rect 237297 66181 237331 66215
rect 222485 63529 222519 63563
rect 216965 56593 216999 56627
rect 237297 56593 237331 56627
rect 238677 66181 238711 66215
rect 385049 66249 385083 66283
rect 240425 62713 240459 62747
rect 238677 56593 238711 56627
rect 239045 57885 239079 57919
rect 210065 48297 210099 48331
rect 218253 56525 218287 56559
rect 180993 46937 181027 46971
rect 218253 46937 218287 46971
rect 222577 54621 222611 54655
rect 158913 46869 158947 46903
rect 182373 46869 182407 46903
rect 158913 29053 158947 29087
rect 163145 38573 163179 38607
rect 182373 37281 182407 37315
rect 210065 46869 210099 46903
rect 221013 46869 221047 46903
rect 210065 37281 210099 37315
rect 219541 38709 219575 38743
rect 207397 37213 207431 37247
rect 163145 28985 163179 29019
rect 181085 34697 181119 34731
rect 181085 28985 181119 29019
rect 182373 31705 182407 31739
rect 182373 28985 182407 29019
rect 183753 27693 183787 27727
rect 158913 27557 158947 27591
rect 156429 19261 156463 19295
rect 158913 19193 158947 19227
rect 181177 27557 181211 27591
rect 239045 48297 239079 48331
rect 222577 45577 222611 45611
rect 237297 46869 237331 46903
rect 221013 37281 221047 37315
rect 237297 37281 237331 37315
rect 238677 46869 238711 46903
rect 238677 37281 238711 37315
rect 239045 38709 239079 38743
rect 239045 37281 239079 37315
rect 385325 38573 385359 38607
rect 219541 35921 219575 35955
rect 385325 28985 385359 29019
rect 207397 27625 207431 27659
rect 226625 28917 226659 28951
rect 183753 26333 183787 26367
rect 216965 27557 216999 27591
rect 181177 17969 181211 18003
rect 183753 26197 183787 26231
rect 207213 22117 207247 22151
rect 183753 16609 183787 16643
rect 200405 19261 200439 19295
rect 156429 12393 156463 12427
rect 183753 13141 183787 13175
rect 183753 8041 183787 8075
rect 185133 12461 185167 12495
rect 207213 17969 207247 18003
rect 200405 9673 200439 9707
rect 216965 9673 216999 9707
rect 219541 27557 219575 27591
rect 239045 28917 239079 28951
rect 226625 19941 226659 19975
rect 237205 27489 237239 27523
rect 222485 19261 222519 19295
rect 222485 11713 222519 11747
rect 219541 9673 219575 9707
rect 237205 9673 237239 9707
rect 238401 27489 238435 27523
rect 239045 22729 239079 22763
rect 257077 19261 257111 19295
rect 257077 12257 257111 12291
rect 385049 19261 385083 19295
rect 238401 9673 238435 9707
rect 385049 9673 385083 9707
rect 185133 4301 185167 4335
rect 222209 5797 222243 5831
rect 93777 4097 93811 4131
rect 84761 4029 84795 4063
rect 42809 3485 42843 3519
rect 42809 3281 42843 3315
rect 84853 4029 84887 4063
rect 84853 3349 84887 3383
rect 84761 3145 84795 3179
rect 220093 3961 220127 3995
rect 170597 3825 170631 3859
rect 167009 3757 167043 3791
rect 162133 3621 162167 3655
rect 162041 3417 162075 3451
rect 162133 3417 162167 3451
rect 162225 3621 162259 3655
rect 167009 3621 167043 3655
rect 211169 3757 211203 3791
rect 170597 3621 170631 3655
rect 174001 3689 174035 3723
rect 174001 3553 174035 3587
rect 201417 3621 201451 3655
rect 93777 3145 93811 3179
rect 107669 3145 107703 3179
rect 111073 3145 111107 3179
rect 111809 3145 111843 3179
rect 111809 3009 111843 3043
rect 111901 3009 111935 3043
rect 121469 2873 121503 2907
rect 121653 2873 121687 2907
rect 107485 2805 107519 2839
rect 202889 3621 202923 3655
rect 202889 3485 202923 3519
rect 206109 3553 206143 3587
rect 201417 1853 201451 1887
rect 220093 3689 220127 3723
rect 220737 3757 220771 3791
rect 211169 3485 211203 3519
rect 220737 3485 220771 3519
rect 230489 4777 230523 4811
rect 226441 3893 226475 3927
rect 224877 3757 224911 3791
rect 229477 3825 229511 3859
rect 229753 3825 229787 3859
rect 224877 3417 224911 3451
rect 226349 3553 226383 3587
rect 226441 3553 226475 3587
rect 222209 3009 222243 3043
rect 234721 4097 234755 4131
rect 234629 3961 234663 3995
rect 234721 3961 234755 3995
rect 234629 3689 234663 3723
rect 306297 3689 306331 3723
rect 275661 3621 275695 3655
rect 304825 3621 304859 3655
rect 230489 3485 230523 3519
rect 233525 3485 233559 3519
rect 226349 3009 226383 3043
rect 243001 3417 243035 3451
rect 306113 3553 306147 3587
rect 306297 3553 306331 3587
rect 275661 3349 275695 3383
rect 243001 3213 243035 3247
rect 233525 3009 233559 3043
rect 319913 3145 319947 3179
rect 325433 3077 325467 3111
rect 319913 2941 319947 2975
rect 320557 3009 320591 3043
rect 320005 2873 320039 2907
rect 325433 2873 325467 2907
rect 206109 1241 206143 1275
rect 255053 2805 255087 2839
rect 255053 561 255087 595
<< metal1 >>
rect 315942 700816 315948 700868
rect 316000 700856 316006 700868
rect 397454 700856 397460 700868
rect 316000 700828 397460 700856
rect 316000 700816 316006 700828
rect 397454 700816 397460 700828
rect 397512 700816 397518 700868
rect 325602 700748 325608 700800
rect 325660 700788 325666 700800
rect 413646 700788 413652 700800
rect 325660 700760 413652 700788
rect 325660 700748 325666 700760
rect 413646 700748 413652 700760
rect 413704 700748 413710 700800
rect 333882 700680 333888 700732
rect 333940 700720 333946 700732
rect 429838 700720 429844 700732
rect 333940 700692 429844 700720
rect 333940 700680 333946 700692
rect 429838 700680 429844 700692
rect 429896 700680 429902 700732
rect 342162 700612 342168 700664
rect 342220 700652 342226 700664
rect 462314 700652 462320 700664
rect 342220 700624 462320 700652
rect 342220 700612 342226 700624
rect 462314 700612 462320 700624
rect 462372 700612 462378 700664
rect 351822 700544 351828 700596
rect 351880 700584 351886 700596
rect 478506 700584 478512 700596
rect 351880 700556 478512 700584
rect 351880 700544 351886 700556
rect 478506 700544 478512 700556
rect 478564 700544 478570 700596
rect 360102 700476 360108 700528
rect 360160 700516 360166 700528
rect 494790 700516 494796 700528
rect 360160 700488 494796 700516
rect 360160 700476 360166 700488
rect 494790 700476 494796 700488
rect 494848 700476 494854 700528
rect 289722 700408 289728 700460
rect 289780 700448 289786 700460
rect 332502 700448 332508 700460
rect 289780 700420 332508 700448
rect 289780 700408 289786 700420
rect 332502 700408 332508 700420
rect 332560 700408 332566 700460
rect 368382 700408 368388 700460
rect 368440 700448 368446 700460
rect 527174 700448 527180 700460
rect 368440 700420 527180 700448
rect 368440 700408 368446 700420
rect 527174 700408 527180 700420
rect 527232 700408 527238 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 273162 700340 273168 700392
rect 273220 700380 273226 700392
rect 283834 700380 283840 700392
rect 273220 700352 283840 700380
rect 273220 700340 273226 700352
rect 283834 700340 283840 700352
rect 283892 700340 283898 700392
rect 299382 700340 299388 700392
rect 299440 700380 299446 700392
rect 348786 700380 348792 700392
rect 299440 700352 348792 700380
rect 299440 700340 299446 700352
rect 348786 700340 348792 700352
rect 348844 700340 348850 700392
rect 376662 700340 376668 700392
rect 376720 700380 376726 700392
rect 543458 700380 543464 700392
rect 376720 700352 543464 700380
rect 376720 700340 376726 700352
rect 543458 700340 543464 700352
rect 543516 700340 543522 700392
rect 281442 700272 281448 700324
rect 281500 700312 281506 700324
rect 300118 700312 300124 700324
rect 281500 700284 300124 700312
rect 281500 700272 281506 700284
rect 300118 700272 300124 700284
rect 300176 700272 300182 700324
rect 307662 700272 307668 700324
rect 307720 700312 307726 700324
rect 364978 700312 364984 700324
rect 307720 700284 364984 700312
rect 307720 700272 307726 700284
rect 364978 700272 364984 700284
rect 365036 700272 365042 700324
rect 386322 700272 386328 700324
rect 386380 700312 386386 700324
rect 559650 700312 559656 700324
rect 386380 700284 559656 700312
rect 386380 700272 386386 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 170306 700204 170312 700256
rect 170364 700244 170370 700256
rect 171042 700244 171048 700256
rect 170364 700216 171048 700244
rect 170364 700204 170370 700216
rect 171042 700204 171048 700216
rect 171100 700204 171106 700256
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 89622 699700 89628 699712
rect 89220 699672 89628 699700
rect 89220 699660 89226 699672
rect 89622 699660 89628 699672
rect 89680 699660 89686 699712
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 264882 699660 264888 699712
rect 264940 699700 264946 699712
rect 267642 699700 267648 699712
rect 264940 699672 267648 699700
rect 264940 699660 264946 699672
rect 267642 699660 267648 699672
rect 267700 699660 267706 699712
rect 8018 698232 8024 698284
rect 8076 698272 8082 698284
rect 8202 698272 8208 698284
rect 8076 698244 8208 698272
rect 8076 698232 8082 698244
rect 8202 698232 8208 698244
rect 8260 698232 8266 698284
rect 137738 698232 137744 698284
rect 137796 698272 137802 698284
rect 137922 698272 137928 698284
rect 137796 698244 137928 698272
rect 137796 698232 137802 698244
rect 137922 698232 137928 698244
rect 137980 698232 137986 698284
rect 393958 696940 393964 696992
rect 394016 696980 394022 696992
rect 580166 696980 580172 696992
rect 394016 696952 580172 696980
rect 394016 696940 394022 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 154114 695512 154120 695564
rect 154172 695552 154178 695564
rect 154206 695552 154212 695564
rect 154172 695524 154212 695552
rect 154172 695512 154178 695524
rect 154206 695512 154212 695524
rect 154264 695512 154270 695564
rect 8113 695487 8171 695493
rect 8113 695453 8125 695487
rect 8159 695484 8171 695487
rect 8202 695484 8208 695496
rect 8159 695456 8208 695484
rect 8159 695453 8171 695456
rect 8113 695447 8171 695453
rect 8202 695444 8208 695456
rect 8260 695444 8266 695496
rect 137833 695487 137891 695493
rect 137833 695453 137845 695487
rect 137879 695484 137891 695487
rect 137922 695484 137928 695496
rect 137879 695456 137928 695484
rect 137879 695453 137891 695456
rect 137833 695447 137891 695453
rect 137922 695444 137928 695456
rect 137980 695444 137986 695496
rect 219069 695487 219127 695493
rect 219069 695453 219081 695487
rect 219115 695484 219127 695487
rect 219158 695484 219164 695496
rect 219115 695456 219164 695484
rect 219115 695453 219127 695456
rect 219069 695447 219127 695453
rect 219158 695444 219164 695456
rect 219216 695444 219222 695496
rect 72513 694127 72571 694133
rect 72513 694093 72525 694127
rect 72559 694124 72571 694127
rect 72694 694124 72700 694136
rect 72559 694096 72700 694124
rect 72559 694093 72571 694096
rect 72513 694087 72571 694093
rect 72694 694084 72700 694096
rect 72752 694084 72758 694136
rect 154206 688576 154212 688628
rect 154264 688616 154270 688628
rect 154390 688616 154396 688628
rect 154264 688588 154396 688616
rect 154264 688576 154270 688588
rect 154390 688576 154396 688588
rect 154448 688576 154454 688628
rect 8110 685896 8116 685908
rect 8071 685868 8116 685896
rect 8110 685856 8116 685868
rect 8168 685856 8174 685908
rect 137830 685896 137836 685908
rect 137791 685868 137836 685896
rect 137830 685856 137836 685868
rect 137888 685856 137894 685908
rect 219066 685896 219072 685908
rect 219027 685868 219072 685896
rect 219066 685856 219072 685868
rect 219124 685856 219130 685908
rect 392578 685856 392584 685908
rect 392636 685896 392642 685908
rect 580166 685896 580172 685908
rect 392636 685868 580172 685896
rect 392636 685856 392642 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 154301 685831 154359 685837
rect 154301 685797 154313 685831
rect 154347 685828 154359 685831
rect 154390 685828 154396 685840
rect 154347 685800 154396 685828
rect 154347 685797 154359 685800
rect 154301 685791 154359 685797
rect 154390 685788 154396 685800
rect 154448 685788 154454 685840
rect 72510 684604 72516 684616
rect 72471 684576 72516 684604
rect 72510 684564 72516 684576
rect 72568 684564 72574 684616
rect 72510 684428 72516 684480
rect 72568 684468 72574 684480
rect 72789 684471 72847 684477
rect 72789 684468 72801 684471
rect 72568 684440 72801 684468
rect 72568 684428 72574 684440
rect 72789 684437 72801 684440
rect 72835 684437 72847 684471
rect 72789 684431 72847 684437
rect 3326 681708 3332 681760
rect 3384 681748 3390 681760
rect 6178 681748 6184 681760
rect 3384 681720 6184 681748
rect 3384 681708 3390 681720
rect 6178 681708 6184 681720
rect 6236 681708 6242 681760
rect 8110 679028 8116 679040
rect 8036 679000 8116 679028
rect 8036 678972 8064 679000
rect 8110 678988 8116 679000
rect 8168 678988 8174 679040
rect 137830 679028 137836 679040
rect 137756 679000 137836 679028
rect 137756 678972 137784 679000
rect 137830 678988 137836 679000
rect 137888 678988 137894 679040
rect 8018 678920 8024 678972
rect 8076 678920 8082 678972
rect 137738 678920 137744 678972
rect 137796 678920 137802 678972
rect 154298 676240 154304 676252
rect 154259 676212 154304 676240
rect 154298 676200 154304 676212
rect 154356 676200 154362 676252
rect 218974 676172 218980 676184
rect 218935 676144 218980 676172
rect 218974 676132 218980 676144
rect 219032 676132 219038 676184
rect 72786 676104 72792 676116
rect 72747 676076 72792 676104
rect 72786 676064 72792 676076
rect 72844 676064 72850 676116
rect 8018 673480 8024 673532
rect 8076 673520 8082 673532
rect 8202 673520 8208 673532
rect 8076 673492 8208 673520
rect 8076 673480 8082 673492
rect 8202 673480 8208 673492
rect 8260 673480 8266 673532
rect 137738 673480 137744 673532
rect 137796 673520 137802 673532
rect 137922 673520 137928 673532
rect 137796 673492 137928 673520
rect 137796 673480 137802 673492
rect 137922 673480 137928 673492
rect 137980 673480 137986 673532
rect 154298 673480 154304 673532
rect 154356 673520 154362 673532
rect 154482 673520 154488 673532
rect 154356 673492 154488 673520
rect 154356 673480 154362 673492
rect 154482 673480 154488 673492
rect 154540 673480 154546 673532
rect 72786 669332 72792 669384
rect 72844 669332 72850 669384
rect 72804 669248 72832 669332
rect 72786 669196 72792 669248
rect 72844 669196 72850 669248
rect 218977 666587 219035 666593
rect 218977 666553 218989 666587
rect 219023 666584 219035 666587
rect 219066 666584 219072 666596
rect 219023 666556 219072 666584
rect 219023 666553 219035 666556
rect 218977 666547 219035 666553
rect 219066 666544 219072 666556
rect 219124 666544 219130 666596
rect 72878 659608 72884 659660
rect 72936 659648 72942 659660
rect 73062 659648 73068 659660
rect 72936 659620 73068 659648
rect 72936 659608 72942 659620
rect 73062 659608 73068 659620
rect 73120 659608 73126 659660
rect 219158 659608 219164 659660
rect 219216 659648 219222 659660
rect 219342 659648 219348 659660
rect 219216 659620 219348 659648
rect 219216 659608 219222 659620
rect 219342 659608 219348 659620
rect 219400 659608 219406 659660
rect 72973 656863 73031 656869
rect 72973 656829 72985 656863
rect 73019 656860 73031 656863
rect 73062 656860 73068 656872
rect 73019 656832 73068 656860
rect 73019 656829 73031 656832
rect 72973 656823 73031 656829
rect 73062 656820 73068 656832
rect 73120 656820 73126 656872
rect 219253 656863 219311 656869
rect 219253 656829 219265 656863
rect 219299 656860 219311 656863
rect 219342 656860 219348 656872
rect 219299 656832 219348 656860
rect 219299 656829 219311 656832
rect 219253 656823 219311 656829
rect 219342 656820 219348 656832
rect 219400 656820 219406 656872
rect 8018 654100 8024 654152
rect 8076 654140 8082 654152
rect 8202 654140 8208 654152
rect 8076 654112 8208 654140
rect 8076 654100 8082 654112
rect 8202 654100 8208 654112
rect 8260 654100 8266 654152
rect 137738 654100 137744 654152
rect 137796 654140 137802 654152
rect 137922 654140 137928 654152
rect 137796 654112 137928 654140
rect 137796 654100 137802 654112
rect 137922 654100 137928 654112
rect 137980 654100 137986 654152
rect 154298 654100 154304 654152
rect 154356 654140 154362 654152
rect 154482 654140 154488 654152
rect 154356 654112 154488 654140
rect 154356 654100 154362 654112
rect 154482 654100 154488 654112
rect 154540 654100 154546 654152
rect 72970 647272 72976 647284
rect 72931 647244 72976 647272
rect 72970 647232 72976 647244
rect 73028 647232 73034 647284
rect 219250 647272 219256 647284
rect 219211 647244 219256 647272
rect 219250 647232 219256 647244
rect 219308 647232 219314 647284
rect 72970 640404 72976 640416
rect 72804 640376 72976 640404
rect 72804 640280 72832 640376
rect 72970 640364 72976 640376
rect 73028 640364 73034 640416
rect 219250 640404 219256 640416
rect 219084 640376 219256 640404
rect 219084 640280 219112 640376
rect 219250 640364 219256 640376
rect 219308 640364 219314 640416
rect 72786 640228 72792 640280
rect 72844 640228 72850 640280
rect 219066 640228 219072 640280
rect 219124 640228 219130 640280
rect 398098 638936 398104 638988
rect 398156 638976 398162 638988
rect 579890 638976 579896 638988
rect 398156 638948 579896 638976
rect 398156 638936 398162 638948
rect 579890 638936 579896 638948
rect 579948 638936 579954 638988
rect 72786 637508 72792 637560
rect 72844 637548 72850 637560
rect 72878 637548 72884 637560
rect 72844 637520 72884 637548
rect 72844 637508 72850 637520
rect 72878 637508 72884 637520
rect 72936 637508 72942 637560
rect 219066 637508 219072 637560
rect 219124 637548 219130 637560
rect 219158 637548 219164 637560
rect 219124 637520 219164 637548
rect 219124 637508 219130 637520
rect 219158 637508 219164 637520
rect 219216 637508 219222 637560
rect 8018 634788 8024 634840
rect 8076 634828 8082 634840
rect 8202 634828 8208 634840
rect 8076 634800 8208 634828
rect 8076 634788 8082 634800
rect 8202 634788 8208 634800
rect 8260 634788 8266 634840
rect 137738 634788 137744 634840
rect 137796 634828 137802 634840
rect 137922 634828 137928 634840
rect 137796 634800 137928 634828
rect 137796 634788 137802 634800
rect 137922 634788 137928 634800
rect 137980 634788 137986 634840
rect 154298 634788 154304 634840
rect 154356 634828 154362 634840
rect 154482 634828 154488 634840
rect 154356 634800 154488 634828
rect 154356 634788 154362 634800
rect 154482 634788 154488 634800
rect 154540 634788 154546 634840
rect 73062 626532 73068 626544
rect 73023 626504 73068 626532
rect 73062 626492 73068 626504
rect 73120 626492 73126 626544
rect 219342 626532 219348 626544
rect 219303 626504 219348 626532
rect 219342 626492 219348 626504
rect 219400 626492 219406 626544
rect 3050 623772 3056 623824
rect 3108 623812 3114 623824
rect 133138 623812 133144 623824
rect 3108 623784 133144 623812
rect 3108 623772 3114 623784
rect 133138 623772 133144 623784
rect 133196 623772 133202 623824
rect 73062 616876 73068 616888
rect 73023 616848 73068 616876
rect 73062 616836 73068 616848
rect 73120 616836 73126 616888
rect 219342 616876 219348 616888
rect 219303 616848 219348 616876
rect 219342 616836 219348 616848
rect 219400 616836 219406 616888
rect 8018 615476 8024 615528
rect 8076 615516 8082 615528
rect 8202 615516 8208 615528
rect 8076 615488 8208 615516
rect 8076 615476 8082 615488
rect 8202 615476 8208 615488
rect 8260 615476 8266 615528
rect 137738 615476 137744 615528
rect 137796 615516 137802 615528
rect 137922 615516 137928 615528
rect 137796 615488 137928 615516
rect 137796 615476 137802 615488
rect 137922 615476 137928 615488
rect 137980 615476 137986 615528
rect 154298 615476 154304 615528
rect 154356 615516 154362 615528
rect 154482 615516 154488 615528
rect 154356 615488 154488 615516
rect 154356 615476 154362 615488
rect 154482 615476 154488 615488
rect 154540 615476 154546 615528
rect 73062 611436 73068 611448
rect 72896 611408 73068 611436
rect 72896 611312 72924 611408
rect 73062 611396 73068 611408
rect 73120 611396 73126 611448
rect 219069 611439 219127 611445
rect 219069 611405 219081 611439
rect 219115 611436 219127 611439
rect 219342 611436 219348 611448
rect 219115 611408 219348 611436
rect 219115 611405 219127 611408
rect 219069 611399 219127 611405
rect 219342 611396 219348 611408
rect 219400 611396 219406 611448
rect 72878 611260 72884 611312
rect 72936 611260 72942 611312
rect 219066 608716 219072 608728
rect 219027 608688 219072 608716
rect 219066 608676 219072 608688
rect 219124 608676 219130 608728
rect 219066 608540 219072 608592
rect 219124 608580 219130 608592
rect 219253 608583 219311 608589
rect 219253 608580 219265 608583
rect 219124 608552 219265 608580
rect 219124 608540 219130 608552
rect 219253 608549 219265 608552
rect 219299 608549 219311 608583
rect 219253 608543 219311 608549
rect 72970 601536 72976 601588
rect 73028 601576 73034 601588
rect 73154 601576 73160 601588
rect 73028 601548 73160 601576
rect 73028 601536 73034 601548
rect 73154 601536 73160 601548
rect 73212 601536 73218 601588
rect 219250 601576 219256 601588
rect 219211 601548 219256 601576
rect 219250 601536 219256 601548
rect 219308 601536 219314 601588
rect 72881 598927 72939 598933
rect 72881 598893 72893 598927
rect 72927 598924 72939 598927
rect 72970 598924 72976 598936
rect 72927 598896 72976 598924
rect 72927 598893 72939 598896
rect 72881 598887 72939 598893
rect 72970 598884 72976 598896
rect 73028 598884 73034 598936
rect 219161 598927 219219 598933
rect 219161 598893 219173 598927
rect 219207 598924 219219 598927
rect 219250 598924 219256 598936
rect 219207 598896 219256 598924
rect 219207 598893 219219 598896
rect 219161 598887 219219 598893
rect 219250 598884 219256 598896
rect 219308 598884 219314 598936
rect 8018 596164 8024 596216
rect 8076 596204 8082 596216
rect 8202 596204 8208 596216
rect 8076 596176 8208 596204
rect 8076 596164 8082 596176
rect 8202 596164 8208 596176
rect 8260 596164 8266 596216
rect 137738 596164 137744 596216
rect 137796 596204 137802 596216
rect 137922 596204 137928 596216
rect 137796 596176 137928 596204
rect 137796 596164 137802 596176
rect 137922 596164 137928 596176
rect 137980 596164 137986 596216
rect 154298 596164 154304 596216
rect 154356 596204 154362 596216
rect 154482 596204 154488 596216
rect 154356 596176 154488 596204
rect 154356 596164 154362 596176
rect 154482 596164 154488 596176
rect 154540 596164 154546 596216
rect 392670 592016 392676 592068
rect 392728 592056 392734 592068
rect 580166 592056 580172 592068
rect 392728 592028 580172 592056
rect 392728 592016 392734 592028
rect 580166 592016 580172 592028
rect 580224 592016 580230 592068
rect 72878 589336 72884 589348
rect 72839 589308 72884 589336
rect 72878 589296 72884 589308
rect 72936 589296 72942 589348
rect 219158 589336 219164 589348
rect 219119 589308 219164 589336
rect 219158 589296 219164 589308
rect 219216 589296 219222 589348
rect 8018 589268 8024 589280
rect 7979 589240 8024 589268
rect 8018 589228 8024 589240
rect 8076 589228 8082 589280
rect 137738 589268 137744 589280
rect 137699 589240 137744 589268
rect 137738 589228 137744 589240
rect 137796 589228 137802 589280
rect 154298 589268 154304 589280
rect 154259 589240 154304 589268
rect 154298 589228 154304 589240
rect 154356 589228 154362 589280
rect 72694 582360 72700 582412
rect 72752 582400 72758 582412
rect 72878 582400 72884 582412
rect 72752 582372 72884 582400
rect 72752 582360 72758 582372
rect 72878 582360 72884 582372
rect 72936 582360 72942 582412
rect 218974 582360 218980 582412
rect 219032 582400 219038 582412
rect 219158 582400 219164 582412
rect 219032 582372 219164 582400
rect 219032 582360 219038 582372
rect 219158 582360 219164 582372
rect 219216 582360 219222 582412
rect 8018 579748 8024 579760
rect 7979 579720 8024 579748
rect 8018 579708 8024 579720
rect 8076 579708 8082 579760
rect 137738 579748 137744 579760
rect 137699 579720 137744 579748
rect 137738 579708 137744 579720
rect 137796 579708 137802 579760
rect 154298 579748 154304 579760
rect 154259 579720 154304 579748
rect 154298 579708 154304 579720
rect 154356 579708 154362 579760
rect 7926 579572 7932 579624
rect 7984 579612 7990 579624
rect 8110 579612 8116 579624
rect 7984 579584 8116 579612
rect 7984 579572 7990 579584
rect 8110 579572 8116 579584
rect 8168 579572 8174 579624
rect 72605 579615 72663 579621
rect 72605 579581 72617 579615
rect 72651 579612 72663 579615
rect 72694 579612 72700 579624
rect 72651 579584 72700 579612
rect 72651 579581 72663 579584
rect 72605 579575 72663 579581
rect 72694 579572 72700 579584
rect 72752 579572 72758 579624
rect 137557 579615 137615 579621
rect 137557 579581 137569 579615
rect 137603 579612 137615 579615
rect 137646 579612 137652 579624
rect 137603 579584 137652 579612
rect 137603 579581 137615 579584
rect 137557 579575 137615 579581
rect 137646 579572 137652 579584
rect 137704 579572 137710 579624
rect 154206 579572 154212 579624
rect 154264 579612 154270 579624
rect 154390 579612 154396 579624
rect 154264 579584 154396 579612
rect 154264 579572 154270 579584
rect 154390 579572 154396 579584
rect 154448 579572 154454 579624
rect 218885 579615 218943 579621
rect 218885 579581 218897 579615
rect 218931 579612 218943 579615
rect 218974 579612 218980 579624
rect 218931 579584 218980 579612
rect 218931 579581 218943 579584
rect 218885 579575 218943 579581
rect 218974 579572 218980 579584
rect 219032 579572 219038 579624
rect 72602 569956 72608 569968
rect 72563 569928 72608 569956
rect 72602 569916 72608 569928
rect 72660 569916 72666 569968
rect 137554 569956 137560 569968
rect 137515 569928 137560 569956
rect 137554 569916 137560 569928
rect 137612 569916 137618 569968
rect 218882 569956 218888 569968
rect 218843 569928 218888 569956
rect 218882 569916 218888 569928
rect 218940 569916 218946 569968
rect 4062 567196 4068 567248
rect 4120 567236 4126 567248
rect 15838 567236 15844 567248
rect 4120 567208 15844 567236
rect 4120 567196 4126 567208
rect 15838 567196 15844 567208
rect 15896 567196 15902 567248
rect 72602 563048 72608 563100
rect 72660 563048 72666 563100
rect 137554 563048 137560 563100
rect 137612 563048 137618 563100
rect 218882 563048 218888 563100
rect 218940 563048 218946 563100
rect 7926 562912 7932 562964
rect 7984 562952 7990 562964
rect 8110 562952 8116 562964
rect 7984 562924 8116 562952
rect 7984 562912 7990 562924
rect 8110 562912 8116 562924
rect 8168 562912 8174 562964
rect 72620 562952 72648 563048
rect 72694 562952 72700 562964
rect 72620 562924 72700 562952
rect 72694 562912 72700 562924
rect 72752 562912 72758 562964
rect 137572 562952 137600 563048
rect 137646 562952 137652 562964
rect 137572 562924 137652 562952
rect 137646 562912 137652 562924
rect 137704 562912 137710 562964
rect 154206 562912 154212 562964
rect 154264 562952 154270 562964
rect 154390 562952 154396 562964
rect 154264 562924 154396 562952
rect 154264 562912 154270 562924
rect 154390 562912 154396 562924
rect 154448 562912 154454 562964
rect 218900 562952 218928 563048
rect 218974 562952 218980 562964
rect 218900 562924 218980 562952
rect 218974 562912 218980 562924
rect 219032 562912 219038 562964
rect 137646 560232 137652 560244
rect 137607 560204 137652 560232
rect 137646 560192 137652 560204
rect 137704 560192 137710 560244
rect 72602 553432 72608 553444
rect 72563 553404 72608 553432
rect 72602 553392 72608 553404
rect 72660 553392 72666 553444
rect 218882 553432 218888 553444
rect 218843 553404 218888 553432
rect 218882 553392 218888 553404
rect 218940 553392 218946 553444
rect 72602 550644 72608 550656
rect 72563 550616 72608 550644
rect 72602 550604 72608 550616
rect 72660 550604 72666 550656
rect 137649 550647 137707 550653
rect 137649 550613 137661 550647
rect 137695 550644 137707 550647
rect 137830 550644 137836 550656
rect 137695 550616 137836 550644
rect 137695 550613 137707 550616
rect 137649 550607 137707 550613
rect 137830 550604 137836 550616
rect 137888 550604 137894 550656
rect 218882 550644 218888 550656
rect 218843 550616 218888 550644
rect 218882 550604 218888 550616
rect 218940 550604 218946 550656
rect 8018 550576 8024 550588
rect 7979 550548 8024 550576
rect 8018 550536 8024 550548
rect 8076 550536 8082 550588
rect 396718 545096 396724 545148
rect 396776 545136 396782 545148
rect 580166 545136 580172 545148
rect 396776 545108 580172 545136
rect 396776 545096 396782 545108
rect 580166 545096 580172 545108
rect 580224 545096 580230 545148
rect 72602 543736 72608 543788
rect 72660 543736 72666 543788
rect 218882 543736 218888 543788
rect 218940 543736 218946 543788
rect 72620 543640 72648 543736
rect 72694 543640 72700 543652
rect 72620 543612 72700 543640
rect 72694 543600 72700 543612
rect 72752 543600 72758 543652
rect 137646 543600 137652 543652
rect 137704 543640 137710 543652
rect 137830 543640 137836 543652
rect 137704 543612 137836 543640
rect 137704 543600 137710 543612
rect 137830 543600 137836 543612
rect 137888 543600 137894 543652
rect 218900 543640 218928 543736
rect 218974 543640 218980 543652
rect 218900 543612 218980 543640
rect 218974 543600 218980 543612
rect 219032 543600 219038 543652
rect 8021 540991 8079 540997
rect 8021 540957 8033 540991
rect 8067 540988 8079 540991
rect 8202 540988 8208 541000
rect 8067 540960 8208 540988
rect 8067 540957 8079 540960
rect 8021 540951 8079 540957
rect 8202 540948 8208 540960
rect 8260 540948 8266 541000
rect 72602 534120 72608 534132
rect 72563 534092 72608 534120
rect 72602 534080 72608 534092
rect 72660 534080 72666 534132
rect 137646 534012 137652 534064
rect 137704 534052 137710 534064
rect 137830 534052 137836 534064
rect 137704 534024 137836 534052
rect 137704 534012 137710 534024
rect 137830 534012 137836 534024
rect 137888 534012 137894 534064
rect 72602 531332 72608 531344
rect 72563 531304 72608 531332
rect 72602 531292 72608 531304
rect 72660 531292 72666 531344
rect 154390 531264 154396 531276
rect 154351 531236 154396 531264
rect 154390 531224 154396 531236
rect 154448 531224 154454 531276
rect 72694 524288 72700 524340
rect 72752 524328 72758 524340
rect 72878 524328 72884 524340
rect 72752 524300 72884 524328
rect 72752 524288 72758 524300
rect 72878 524288 72884 524300
rect 72936 524288 72942 524340
rect 218974 524288 218980 524340
rect 219032 524328 219038 524340
rect 219158 524328 219164 524340
rect 219032 524300 219164 524328
rect 219032 524288 219038 524300
rect 219158 524288 219164 524300
rect 219216 524288 219222 524340
rect 8202 521636 8208 521688
rect 8260 521676 8266 521688
rect 8386 521676 8392 521688
rect 8260 521648 8392 521676
rect 8260 521636 8266 521648
rect 8386 521636 8392 521648
rect 8444 521636 8450 521688
rect 137922 521636 137928 521688
rect 137980 521676 137986 521688
rect 138106 521676 138112 521688
rect 137980 521648 138112 521676
rect 137980 521636 137986 521648
rect 138106 521636 138112 521648
rect 138164 521636 138170 521688
rect 154393 521679 154451 521685
rect 154393 521645 154405 521679
rect 154439 521676 154451 521679
rect 154482 521676 154488 521688
rect 154439 521648 154488 521676
rect 154439 521645 154451 521648
rect 154393 521639 154451 521645
rect 154482 521636 154488 521648
rect 154540 521636 154546 521688
rect 154390 511952 154396 511964
rect 154351 511924 154396 511952
rect 154390 511912 154396 511924
rect 154448 511912 154454 511964
rect 3326 509736 3332 509788
rect 3384 509776 3390 509788
rect 10318 509776 10324 509788
rect 3384 509748 10324 509776
rect 3384 509736 3390 509748
rect 10318 509736 10324 509748
rect 10376 509736 10382 509788
rect 8202 502324 8208 502376
rect 8260 502364 8266 502376
rect 8386 502364 8392 502376
rect 8260 502336 8392 502364
rect 8260 502324 8266 502336
rect 8386 502324 8392 502336
rect 8444 502324 8450 502376
rect 72602 502324 72608 502376
rect 72660 502364 72666 502376
rect 73062 502364 73068 502376
rect 72660 502336 73068 502364
rect 72660 502324 72666 502336
rect 73062 502324 73068 502336
rect 73120 502324 73126 502376
rect 137922 502324 137928 502376
rect 137980 502364 137986 502376
rect 138106 502364 138112 502376
rect 137980 502336 138112 502364
rect 137980 502324 137986 502336
rect 138106 502324 138112 502336
rect 138164 502324 138170 502376
rect 154393 502367 154451 502373
rect 154393 502333 154405 502367
rect 154439 502364 154451 502367
rect 154482 502364 154488 502376
rect 154439 502336 154488 502364
rect 154439 502333 154451 502336
rect 154393 502327 154451 502333
rect 154482 502324 154488 502336
rect 154540 502324 154546 502376
rect 218882 502324 218888 502376
rect 218940 502364 218946 502376
rect 219342 502364 219348 502376
rect 218940 502336 219348 502364
rect 218940 502324 218946 502336
rect 219342 502324 219348 502336
rect 219400 502324 219406 502376
rect 392762 498176 392768 498228
rect 392820 498216 392826 498228
rect 579982 498216 579988 498228
rect 392820 498188 579988 498216
rect 392820 498176 392826 498188
rect 579982 498176 579988 498188
rect 580040 498176 580046 498228
rect 137646 492600 137652 492652
rect 137704 492640 137710 492652
rect 137830 492640 137836 492652
rect 137704 492612 137836 492640
rect 137704 492600 137710 492612
rect 137830 492600 137836 492612
rect 137888 492600 137894 492652
rect 154206 492600 154212 492652
rect 154264 492640 154270 492652
rect 154390 492640 154396 492652
rect 154264 492612 154396 492640
rect 154264 492600 154270 492612
rect 154390 492600 154396 492612
rect 154448 492600 154454 492652
rect 8110 485800 8116 485852
rect 8168 485800 8174 485852
rect 400858 485800 400864 485852
rect 400916 485840 400922 485852
rect 579982 485840 579988 485852
rect 400916 485812 579988 485840
rect 400916 485800 400922 485812
rect 579982 485800 579988 485812
rect 580040 485800 580046 485852
rect 8128 485772 8156 485800
rect 8202 485772 8208 485784
rect 8128 485744 8208 485772
rect 8202 485732 8208 485744
rect 8260 485732 8266 485784
rect 7926 482944 7932 482996
rect 7984 482984 7990 482996
rect 8202 482984 8208 482996
rect 7984 482956 8208 482984
rect 7984 482944 7990 482956
rect 8202 482944 8208 482956
rect 8260 482944 8266 482996
rect 72878 480224 72884 480276
rect 72936 480264 72942 480276
rect 73062 480264 73068 480276
rect 72936 480236 73068 480264
rect 72936 480224 72942 480236
rect 73062 480224 73068 480236
rect 73120 480224 73126 480276
rect 219158 480224 219164 480276
rect 219216 480264 219222 480276
rect 219342 480264 219348 480276
rect 219216 480236 219348 480264
rect 219216 480224 219222 480236
rect 219342 480224 219348 480236
rect 219400 480224 219406 480276
rect 137738 466528 137744 466540
rect 137664 466500 137744 466528
rect 8110 466420 8116 466472
rect 8168 466420 8174 466472
rect 8128 466392 8156 466420
rect 137664 466404 137692 466500
rect 137738 466488 137744 466500
rect 137796 466488 137802 466540
rect 154298 466420 154304 466472
rect 154356 466460 154362 466472
rect 154482 466460 154488 466472
rect 154356 466432 154488 466460
rect 154356 466420 154362 466432
rect 154482 466420 154488 466432
rect 154540 466420 154546 466472
rect 8202 466392 8208 466404
rect 8128 466364 8208 466392
rect 8202 466352 8208 466364
rect 8260 466352 8266 466404
rect 137646 466352 137652 466404
rect 137704 466352 137710 466404
rect 137370 463632 137376 463684
rect 137428 463672 137434 463684
rect 137646 463672 137652 463684
rect 137428 463644 137652 463672
rect 137428 463632 137434 463644
rect 137646 463632 137652 463644
rect 137704 463632 137710 463684
rect 395338 462340 395344 462392
rect 395396 462380 395402 462392
rect 579982 462380 579988 462392
rect 395396 462352 579988 462380
rect 395396 462340 395402 462352
rect 579982 462340 579988 462352
rect 580040 462340 580046 462392
rect 72878 460912 72884 460964
rect 72936 460952 72942 460964
rect 73062 460952 73068 460964
rect 72936 460924 73068 460952
rect 72936 460912 72942 460924
rect 73062 460912 73068 460924
rect 73120 460912 73126 460964
rect 219158 460912 219164 460964
rect 219216 460952 219222 460964
rect 219342 460952 219348 460964
rect 219216 460924 219348 460952
rect 219216 460912 219222 460924
rect 219342 460912 219348 460924
rect 219400 460912 219406 460964
rect 7929 454019 7987 454025
rect 7929 453985 7941 454019
rect 7975 454016 7987 454019
rect 8018 454016 8024 454028
rect 7975 453988 8024 454016
rect 7975 453985 7987 453988
rect 7929 453979 7987 453985
rect 8018 453976 8024 453988
rect 8076 453976 8082 454028
rect 154209 454019 154267 454025
rect 154209 453985 154221 454019
rect 154255 454016 154267 454019
rect 154298 454016 154304 454028
rect 154255 453988 154304 454016
rect 154255 453985 154267 453988
rect 154209 453979 154267 453985
rect 154298 453976 154304 453988
rect 154356 453976 154362 454028
rect 3326 451392 3332 451444
rect 3384 451432 3390 451444
rect 11698 451432 11704 451444
rect 3384 451404 11704 451432
rect 3384 451392 3390 451404
rect 11698 451392 11704 451404
rect 11756 451392 11762 451444
rect 399478 451256 399484 451308
rect 399536 451296 399542 451308
rect 579982 451296 579988 451308
rect 399536 451268 579988 451296
rect 399536 451256 399542 451268
rect 579982 451256 579988 451268
rect 580040 451256 580046 451308
rect 137554 447108 137560 447160
rect 137612 447108 137618 447160
rect 137572 447080 137600 447108
rect 137646 447080 137652 447092
rect 137572 447052 137652 447080
rect 137646 447040 137652 447052
rect 137704 447040 137710 447092
rect 7926 444428 7932 444440
rect 7887 444400 7932 444428
rect 7926 444388 7932 444400
rect 7984 444388 7990 444440
rect 154206 444428 154212 444440
rect 154167 444400 154212 444428
rect 154206 444388 154212 444400
rect 154264 444388 154270 444440
rect 72970 444320 72976 444372
rect 73028 444360 73034 444372
rect 73154 444360 73160 444372
rect 73028 444332 73160 444360
rect 73028 444320 73034 444332
rect 73154 444320 73160 444332
rect 73212 444320 73218 444372
rect 219250 444320 219256 444372
rect 219308 444360 219314 444372
rect 219434 444360 219440 444372
rect 219308 444332 219440 444360
rect 219308 444320 219314 444332
rect 219434 444320 219440 444332
rect 219492 444320 219498 444372
rect 3326 437656 3332 437708
rect 3384 437696 3390 437708
rect 4798 437696 4804 437708
rect 3384 437668 4804 437696
rect 3384 437656 3390 437668
rect 4798 437656 4804 437668
rect 4856 437656 4862 437708
rect 8018 427796 8024 427848
rect 8076 427796 8082 427848
rect 137738 427796 137744 427848
rect 137796 427796 137802 427848
rect 154298 427796 154304 427848
rect 154356 427796 154362 427848
rect 8036 427768 8064 427796
rect 8110 427768 8116 427780
rect 8036 427740 8116 427768
rect 8110 427728 8116 427740
rect 8168 427728 8174 427780
rect 137756 427768 137784 427796
rect 137830 427768 137836 427780
rect 137756 427740 137836 427768
rect 137830 427728 137836 427740
rect 137888 427728 137894 427780
rect 154316 427768 154344 427796
rect 154390 427768 154396 427780
rect 154316 427740 154396 427768
rect 154390 427728 154396 427740
rect 154448 427728 154454 427780
rect 7834 425008 7840 425060
rect 7892 425048 7898 425060
rect 8110 425048 8116 425060
rect 7892 425020 8116 425048
rect 7892 425008 7898 425020
rect 8110 425008 8116 425020
rect 8168 425008 8174 425060
rect 137554 425008 137560 425060
rect 137612 425048 137618 425060
rect 137830 425048 137836 425060
rect 137612 425020 137836 425048
rect 137612 425008 137618 425020
rect 137830 425008 137836 425020
rect 137888 425008 137894 425060
rect 154114 425008 154120 425060
rect 154172 425048 154178 425060
rect 154390 425048 154396 425060
rect 154172 425020 154396 425048
rect 154172 425008 154178 425020
rect 154390 425008 154396 425020
rect 154448 425008 154454 425060
rect 72694 418248 72700 418260
rect 72620 418220 72700 418248
rect 72620 418124 72648 418220
rect 72694 418208 72700 418220
rect 72752 418208 72758 418260
rect 218974 418248 218980 418260
rect 218900 418220 218980 418248
rect 218900 418124 218928 418220
rect 218974 418208 218980 418220
rect 219032 418208 219038 418260
rect 72602 418072 72608 418124
rect 72660 418072 72666 418124
rect 218882 418072 218888 418124
rect 218940 418072 218946 418124
rect 392854 415420 392860 415472
rect 392912 415460 392918 415472
rect 580074 415460 580080 415472
rect 392912 415432 580080 415460
rect 392912 415420 392918 415432
rect 580074 415420 580080 415432
rect 580132 415420 580138 415472
rect 263594 415352 263600 415404
rect 263652 415392 263658 415404
rect 264882 415392 264888 415404
rect 263652 415364 264888 415392
rect 263652 415352 263658 415364
rect 264882 415352 264888 415364
rect 264940 415352 264946 415404
rect 298370 415352 298376 415404
rect 298428 415392 298434 415404
rect 299382 415392 299388 415404
rect 298428 415364 299388 415392
rect 298428 415352 298434 415364
rect 299382 415352 299388 415364
rect 299440 415352 299446 415404
rect 359274 415352 359280 415404
rect 359332 415392 359338 415404
rect 360102 415392 360108 415404
rect 359332 415364 360108 415392
rect 359332 415352 359338 415364
rect 360102 415352 360108 415364
rect 360160 415352 360166 415404
rect 385310 415352 385316 415404
rect 385368 415392 385374 415404
rect 386322 415392 386328 415404
rect 385368 415364 386328 415392
rect 385368 415352 385374 415364
rect 386322 415352 386328 415364
rect 386380 415352 386386 415404
rect 154298 415148 154304 415200
rect 154356 415188 154362 415200
rect 220170 415188 220176 415200
rect 154356 415160 220176 415188
rect 154356 415148 154362 415160
rect 220170 415148 220176 415160
rect 220228 415148 220234 415200
rect 137738 415080 137744 415132
rect 137796 415120 137802 415132
rect 211430 415120 211436 415132
rect 137796 415092 211436 415120
rect 137796 415080 137802 415092
rect 211430 415080 211436 415092
rect 211488 415080 211494 415132
rect 350534 415080 350540 415132
rect 350592 415120 350598 415132
rect 351822 415120 351828 415132
rect 350592 415092 351828 415120
rect 350592 415080 350598 415092
rect 351822 415080 351828 415092
rect 351880 415080 351886 415132
rect 106182 415012 106188 415064
rect 106240 415052 106246 415064
rect 202414 415052 202420 415064
rect 106240 415024 202420 415052
rect 106240 415012 106246 415024
rect 202414 415012 202420 415024
rect 202472 415012 202478 415064
rect 89622 414944 89628 414996
rect 89680 414984 89686 414996
rect 194042 414984 194048 414996
rect 89680 414956 194048 414984
rect 89680 414944 89686 414956
rect 194042 414944 194048 414956
rect 194100 414944 194106 414996
rect 72602 414876 72608 414928
rect 72660 414916 72666 414928
rect 185394 414916 185400 414928
rect 72660 414888 185400 414916
rect 72660 414876 72666 414888
rect 185394 414876 185400 414888
rect 185452 414876 185458 414928
rect 41322 414808 41328 414860
rect 41380 414848 41386 414860
rect 176654 414848 176660 414860
rect 41380 414820 176660 414848
rect 41380 414808 41386 414820
rect 176654 414808 176660 414820
rect 176712 414808 176718 414860
rect 218882 414808 218888 414860
rect 218940 414848 218946 414860
rect 246206 414848 246212 414860
rect 218940 414820 246212 414848
rect 218940 414808 218946 414820
rect 246206 414808 246212 414820
rect 246264 414808 246270 414860
rect 24762 414740 24768 414792
rect 24820 414780 24826 414792
rect 168006 414780 168012 414792
rect 24820 414752 168012 414780
rect 24820 414740 24826 414752
rect 168006 414740 168012 414752
rect 168064 414740 168070 414792
rect 202782 414740 202788 414792
rect 202840 414780 202846 414792
rect 237558 414780 237564 414792
rect 202840 414752 237564 414780
rect 202840 414740 202846 414752
rect 237558 414740 237564 414752
rect 237616 414740 237622 414792
rect 8018 414672 8024 414724
rect 8076 414712 8082 414724
rect 159358 414712 159364 414724
rect 8076 414684 159364 414712
rect 8076 414672 8082 414684
rect 159358 414672 159364 414684
rect 159416 414672 159422 414724
rect 171042 414672 171048 414724
rect 171100 414712 171106 414724
rect 228818 414712 228824 414724
rect 171100 414684 228824 414712
rect 171100 414672 171106 414684
rect 228818 414672 228824 414684
rect 228876 414672 228882 414724
rect 235902 414672 235908 414724
rect 235960 414712 235966 414724
rect 254946 414712 254952 414724
rect 235960 414684 254952 414712
rect 235960 414672 235966 414684
rect 254946 414672 254952 414684
rect 255004 414672 255010 414724
rect 272334 414672 272340 414724
rect 272392 414712 272398 414724
rect 273162 414712 273168 414724
rect 272392 414684 273168 414712
rect 272392 414672 272398 414684
rect 273162 414672 273168 414684
rect 273220 414672 273226 414724
rect 324498 414196 324504 414248
rect 324556 414236 324562 414248
rect 325602 414236 325608 414248
rect 324556 414208 325608 414236
rect 324556 414196 324562 414208
rect 325602 414196 325608 414208
rect 325660 414196 325666 414248
rect 579890 412564 579896 412616
rect 579948 412604 579954 412616
rect 580258 412604 580264 412616
rect 579948 412576 580264 412604
rect 579948 412564 579954 412576
rect 580258 412564 580264 412576
rect 580316 412564 580322 412616
rect 3510 409776 3516 409828
rect 3568 409816 3574 409828
rect 151814 409816 151820 409828
rect 3568 409788 151820 409816
rect 3568 409776 3574 409788
rect 151814 409776 151820 409788
rect 151872 409776 151878 409828
rect 391934 409232 391940 409284
rect 391992 409272 391998 409284
rect 393958 409272 393964 409284
rect 391992 409244 393964 409272
rect 391992 409232 391998 409244
rect 393958 409232 393964 409244
rect 394016 409232 394022 409284
rect 393958 404336 393964 404388
rect 394016 404376 394022 404388
rect 580074 404376 580080 404388
rect 394016 404348 580080 404376
rect 394016 404336 394022 404348
rect 580074 404336 580080 404348
rect 580132 404336 580138 404388
rect 3418 404268 3424 404320
rect 3476 404308 3482 404320
rect 152366 404308 152372 404320
rect 3476 404280 152372 404308
rect 3476 404268 3482 404280
rect 152366 404268 152372 404280
rect 152424 404268 152430 404320
rect 6178 398760 6184 398812
rect 6236 398800 6242 398812
rect 153102 398800 153108 398812
rect 6236 398772 153108 398800
rect 6236 398760 6242 398772
rect 153102 398760 153108 398772
rect 153160 398760 153166 398812
rect 391934 398760 391940 398812
rect 391992 398800 391998 398812
rect 580074 398800 580080 398812
rect 391992 398772 580080 398800
rect 391992 398760 391998 398772
rect 580074 398760 580080 398772
rect 580132 398760 580138 398812
rect 391934 394612 391940 394664
rect 391992 394652 391998 394664
rect 580350 394652 580356 394664
rect 391992 394624 580356 394652
rect 391992 394612 391998 394624
rect 580350 394612 580356 394624
rect 580408 394612 580414 394664
rect 3694 393252 3700 393304
rect 3752 393292 3758 393304
rect 153102 393292 153108 393304
rect 3752 393264 153108 393292
rect 3752 393252 3758 393264
rect 153102 393252 153108 393264
rect 153160 393252 153166 393304
rect 391934 389104 391940 389156
rect 391992 389144 391998 389156
rect 398098 389144 398104 389156
rect 391992 389116 398104 389144
rect 391992 389104 391998 389116
rect 398098 389104 398104 389116
rect 398156 389104 398162 389156
rect 3602 386316 3608 386368
rect 3660 386356 3666 386368
rect 153102 386356 153108 386368
rect 3660 386328 153108 386356
rect 3660 386316 3666 386328
rect 153102 386316 153108 386328
rect 153160 386316 153166 386368
rect 391934 383596 391940 383648
rect 391992 383636 391998 383648
rect 580442 383636 580448 383648
rect 391992 383608 580448 383636
rect 391992 383596 391998 383608
rect 580442 383596 580448 383608
rect 580500 383596 580506 383648
rect 133138 380808 133144 380860
rect 133196 380848 133202 380860
rect 152550 380848 152556 380860
rect 133196 380820 152556 380848
rect 133196 380808 133202 380820
rect 152550 380808 152556 380820
rect 152608 380808 152614 380860
rect 391934 378088 391940 378140
rect 391992 378128 391998 378140
rect 580534 378128 580540 378140
rect 391992 378100 580540 378128
rect 391992 378088 391998 378100
rect 580534 378088 580540 378100
rect 580592 378088 580598 378140
rect 3878 375300 3884 375352
rect 3936 375340 3942 375352
rect 152550 375340 152556 375352
rect 3936 375312 152556 375340
rect 3936 375300 3942 375312
rect 152550 375300 152556 375312
rect 152608 375300 152614 375352
rect 3786 369792 3792 369844
rect 3844 369832 3850 369844
rect 152918 369832 152924 369844
rect 3844 369804 152924 369832
rect 3844 369792 3850 369804
rect 152918 369792 152924 369804
rect 152976 369792 152982 369844
rect 392578 368500 392584 368552
rect 392636 368540 392642 368552
rect 580074 368540 580080 368552
rect 392636 368512 580080 368540
rect 392636 368500 392642 368512
rect 580074 368500 580080 368512
rect 580132 368500 580138 368552
rect 391934 367004 391940 367056
rect 391992 367044 391998 367056
rect 580626 367044 580632 367056
rect 391992 367016 580632 367044
rect 391992 367004 391998 367016
rect 580626 367004 580632 367016
rect 580684 367004 580690 367056
rect 15838 364284 15844 364336
rect 15896 364324 15902 364336
rect 153102 364324 153108 364336
rect 15896 364296 153108 364324
rect 15896 364284 15902 364296
rect 153102 364284 153108 364296
rect 153160 364284 153166 364336
rect 391934 362856 391940 362908
rect 391992 362896 391998 362908
rect 580718 362896 580724 362908
rect 391992 362868 580724 362896
rect 391992 362856 391998 362868
rect 580718 362856 580724 362868
rect 580776 362856 580782 362908
rect 4062 358708 4068 358760
rect 4120 358748 4126 358760
rect 153102 358748 153108 358760
rect 4120 358720 153108 358748
rect 4120 358708 4126 358720
rect 153102 358708 153108 358720
rect 153160 358708 153166 358760
rect 392670 357416 392676 357468
rect 392728 357456 392734 357468
rect 580074 357456 580080 357468
rect 392728 357428 580080 357456
rect 392728 357416 392734 357428
rect 580074 357416 580080 357428
rect 580132 357416 580138 357468
rect 391934 357348 391940 357400
rect 391992 357388 391998 357400
rect 396718 357388 396724 357400
rect 391992 357360 396724 357388
rect 391992 357348 391998 357360
rect 396718 357348 396724 357360
rect 396776 357348 396782 357400
rect 3970 353200 3976 353252
rect 4028 353240 4034 353252
rect 153102 353240 153108 353252
rect 4028 353212 153108 353240
rect 4028 353200 4034 353212
rect 153102 353200 153108 353212
rect 153160 353200 153166 353252
rect 391934 351840 391940 351892
rect 391992 351880 391998 351892
rect 580810 351880 580816 351892
rect 391992 351852 580816 351880
rect 391992 351840 391998 351852
rect 580810 351840 580816 351852
rect 580868 351840 580874 351892
rect 10318 347692 10324 347744
rect 10376 347732 10382 347744
rect 152918 347732 152924 347744
rect 10376 347704 152924 347732
rect 10376 347692 10382 347704
rect 152918 347692 152924 347704
rect 152976 347692 152982 347744
rect 391934 346332 391940 346384
rect 391992 346372 391998 346384
rect 580902 346372 580908 346384
rect 391992 346344 580908 346372
rect 391992 346332 391998 346344
rect 580902 346332 580908 346344
rect 580960 346332 580966 346384
rect 3326 342184 3332 342236
rect 3384 342224 3390 342236
rect 152550 342224 152556 342236
rect 3384 342196 152556 342224
rect 3384 342184 3390 342196
rect 152550 342184 152556 342196
rect 152608 342184 152614 342236
rect 4798 336676 4804 336728
rect 4856 336716 4862 336728
rect 153102 336716 153108 336728
rect 4856 336688 153108 336716
rect 4856 336676 4862 336688
rect 153102 336676 153108 336688
rect 153160 336676 153166 336728
rect 391934 336676 391940 336728
rect 391992 336716 391998 336728
rect 400858 336716 400864 336728
rect 391992 336688 400864 336716
rect 391992 336676 391998 336688
rect 400858 336676 400864 336688
rect 400916 336676 400922 336728
rect 11698 331168 11704 331220
rect 11756 331208 11762 331220
rect 153102 331208 153108 331220
rect 11756 331180 153108 331208
rect 11756 331168 11762 331180
rect 153102 331168 153108 331180
rect 153160 331168 153166 331220
rect 391934 330352 391940 330404
rect 391992 330392 391998 330404
rect 395338 330392 395344 330404
rect 391992 330364 395344 330392
rect 391992 330352 391998 330364
rect 395338 330352 395344 330364
rect 395396 330352 395402 330404
rect 391934 325592 391940 325644
rect 391992 325632 391998 325644
rect 399478 325632 399484 325644
rect 391992 325604 399484 325632
rect 391992 325592 391998 325604
rect 399478 325592 399484 325604
rect 399536 325592 399542 325644
rect 3602 324232 3608 324284
rect 3660 324272 3666 324284
rect 153102 324272 153108 324284
rect 3660 324244 153108 324272
rect 3660 324232 3666 324244
rect 153102 324232 153108 324244
rect 153160 324232 153166 324284
rect 579890 322736 579896 322788
rect 579948 322776 579954 322788
rect 580166 322776 580172 322788
rect 579948 322748 580172 322776
rect 579948 322736 579954 322748
rect 580166 322736 580172 322748
rect 580224 322736 580230 322788
rect 392762 321580 392768 321632
rect 392820 321620 392826 321632
rect 580166 321620 580172 321632
rect 392820 321592 580172 321620
rect 392820 321580 392826 321592
rect 580166 321580 580172 321592
rect 580224 321580 580230 321632
rect 391934 320084 391940 320136
rect 391992 320124 391998 320136
rect 579890 320124 579896 320136
rect 391992 320096 579896 320124
rect 391992 320084 391998 320096
rect 579890 320084 579896 320096
rect 579948 320084 579954 320136
rect 3510 318724 3516 318776
rect 3568 318764 3574 318776
rect 153102 318764 153108 318776
rect 3568 318736 153108 318764
rect 3568 318724 3574 318736
rect 153102 318724 153108 318736
rect 153160 318724 153166 318776
rect 3418 313216 3424 313268
rect 3476 313256 3482 313268
rect 152366 313256 152372 313268
rect 3476 313228 152372 313256
rect 3476 313216 3482 313228
rect 152366 313216 152372 313228
rect 152424 313216 152430 313268
rect 392854 310496 392860 310548
rect 392912 310536 392918 310548
rect 579614 310536 579620 310548
rect 392912 310508 579620 310536
rect 392912 310496 392918 310508
rect 579614 310496 579620 310508
rect 579672 310496 579678 310548
rect 391934 309544 391940 309596
rect 391992 309584 391998 309596
rect 393958 309584 393964 309596
rect 391992 309556 393964 309584
rect 391992 309544 391998 309556
rect 393958 309544 393964 309556
rect 394016 309544 394022 309596
rect 3050 307708 3056 307760
rect 3108 307748 3114 307760
rect 152550 307748 152556 307760
rect 3108 307720 152556 307748
rect 3108 307708 3114 307720
rect 152550 307708 152556 307720
rect 152608 307708 152614 307760
rect 391934 304920 391940 304972
rect 391992 304960 391998 304972
rect 580258 304960 580264 304972
rect 391992 304932 580264 304960
rect 391992 304920 391998 304932
rect 580258 304920 580264 304932
rect 580316 304920 580322 304972
rect 3786 302132 3792 302184
rect 3844 302172 3850 302184
rect 153102 302172 153108 302184
rect 3844 302144 153108 302172
rect 3844 302132 3850 302144
rect 153102 302132 153108 302144
rect 153160 302132 153166 302184
rect 3694 296624 3700 296676
rect 3752 296664 3758 296676
rect 152734 296664 152740 296676
rect 3752 296636 152740 296664
rect 3752 296624 3758 296636
rect 152734 296624 152740 296636
rect 152792 296624 152798 296676
rect 3418 289824 3424 289876
rect 3476 289864 3482 289876
rect 152182 289864 152188 289876
rect 3476 289836 152188 289864
rect 3476 289824 3482 289836
rect 152182 289824 152188 289836
rect 152240 289824 152246 289876
rect 391934 288328 391940 288380
rect 391992 288368 391998 288380
rect 580350 288368 580356 288380
rect 391992 288340 580356 288368
rect 391992 288328 391998 288340
rect 580350 288328 580356 288340
rect 580408 288328 580414 288380
rect 2958 284316 2964 284368
rect 3016 284356 3022 284368
rect 151998 284356 152004 284368
rect 3016 284328 152004 284356
rect 3016 284316 3022 284328
rect 151998 284316 152004 284328
rect 152056 284316 152062 284368
rect 3510 280100 3516 280152
rect 3568 280140 3574 280152
rect 152918 280140 152924 280152
rect 3568 280112 152924 280140
rect 3568 280100 3574 280112
rect 152918 280100 152924 280112
rect 152976 280100 152982 280152
rect 392578 274660 392584 274712
rect 392636 274700 392642 274712
rect 580166 274700 580172 274712
rect 392636 274672 580172 274700
rect 392636 274660 392642 274672
rect 580166 274660 580172 274672
rect 580224 274660 580230 274712
rect 391934 273164 391940 273216
rect 391992 273204 391998 273216
rect 580258 273204 580264 273216
rect 391992 273176 580264 273204
rect 391992 273164 391998 273176
rect 580258 273164 580264 273176
rect 580316 273164 580322 273216
rect 3510 267724 3516 267776
rect 3568 267764 3574 267776
rect 153102 267764 153108 267776
rect 3568 267736 153108 267764
rect 3568 267724 3574 267736
rect 153102 267724 153108 267736
rect 153160 267724 153166 267776
rect 391934 263576 391940 263628
rect 391992 263616 391998 263628
rect 579798 263616 579804 263628
rect 391992 263588 579804 263616
rect 391992 263576 391998 263588
rect 579798 263576 579804 263588
rect 579856 263576 579862 263628
rect 3418 262216 3424 262268
rect 3476 262256 3482 262268
rect 153102 262256 153108 262268
rect 3476 262228 153108 262256
rect 3476 262216 3482 262228
rect 153102 262216 153108 262228
rect 153160 262216 153166 262268
rect 391934 252492 391940 252544
rect 391992 252532 391998 252544
rect 579798 252532 579804 252544
rect 391992 252504 579804 252532
rect 391992 252492 391998 252504
rect 579798 252492 579804 252504
rect 579856 252492 579862 252544
rect 3418 249772 3424 249824
rect 3476 249812 3482 249824
rect 153102 249812 153108 249824
rect 3476 249784 153108 249812
rect 3476 249772 3482 249784
rect 153102 249772 153108 249784
rect 153160 249772 153166 249824
rect 3694 233248 3700 233300
rect 3752 233288 3758 233300
rect 153102 233288 153108 233300
rect 3752 233260 153108 233288
rect 3752 233248 3758 233260
rect 153102 233248 153108 233260
rect 153160 233248 153166 233300
rect 392762 229032 392768 229084
rect 392820 229072 392826 229084
rect 580166 229072 580172 229084
rect 392820 229044 580172 229072
rect 392820 229032 392826 229044
rect 580166 229032 580172 229044
rect 580224 229032 580230 229084
rect 3510 223524 3516 223576
rect 3568 223564 3574 223576
rect 152458 223564 152464 223576
rect 3568 223536 152464 223564
rect 3568 223524 3574 223536
rect 152458 223524 152464 223536
rect 152516 223524 152522 223576
rect 392670 217948 392676 218000
rect 392728 217988 392734 218000
rect 580166 217988 580172 218000
rect 392728 217960 580172 217988
rect 392728 217948 392734 217960
rect 580166 217948 580172 217960
rect 580224 217948 580230 218000
rect 3602 216656 3608 216708
rect 3660 216696 3666 216708
rect 153010 216696 153016 216708
rect 3660 216668 153016 216696
rect 3660 216656 3666 216668
rect 153010 216656 153016 216668
rect 153068 216656 153074 216708
rect 391934 208360 391940 208412
rect 391992 208400 391998 208412
rect 395338 208400 395344 208412
rect 391992 208372 395344 208400
rect 391992 208360 391998 208372
rect 395338 208360 395344 208372
rect 395396 208360 395402 208412
rect 3142 208292 3148 208344
rect 3200 208332 3206 208344
rect 152550 208332 152556 208344
rect 3200 208304 152556 208332
rect 3200 208292 3206 208304
rect 152550 208292 152556 208304
rect 152608 208292 152614 208344
rect 392578 205572 392584 205624
rect 392636 205612 392642 205624
rect 579798 205612 579804 205624
rect 392636 205584 579804 205612
rect 392636 205572 392642 205584
rect 579798 205572 579804 205584
rect 579856 205572 579862 205624
rect 3510 200132 3516 200184
rect 3568 200172 3574 200184
rect 151998 200172 152004 200184
rect 3568 200144 152004 200172
rect 3568 200132 3574 200144
rect 151998 200132 152004 200144
rect 152056 200132 152062 200184
rect 3418 182180 3424 182232
rect 3476 182220 3482 182232
rect 152458 182220 152464 182232
rect 3476 182192 152464 182220
rect 3476 182180 3482 182192
rect 152458 182180 152464 182192
rect 152516 182180 152522 182232
rect 392486 182112 392492 182164
rect 392544 182152 392550 182164
rect 580166 182152 580172 182164
rect 392544 182124 580172 182152
rect 392544 182112 392550 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 3050 180752 3056 180804
rect 3108 180792 3114 180804
rect 152642 180792 152648 180804
rect 3108 180764 152648 180792
rect 3108 180752 3114 180764
rect 152642 180752 152648 180764
rect 152700 180752 152706 180804
rect 391934 176672 391940 176724
rect 391992 176712 391998 176724
rect 519078 176712 519084 176724
rect 391992 176684 519084 176712
rect 391992 176672 391998 176684
rect 519078 176672 519084 176684
rect 519136 176672 519142 176724
rect 188062 173992 188068 174004
rect 188023 173964 188068 173992
rect 188062 173952 188068 173964
rect 188120 173952 188126 174004
rect 211062 173816 211068 173868
rect 211120 173856 211126 173868
rect 220081 173859 220139 173865
rect 220081 173856 220093 173859
rect 211120 173828 220093 173856
rect 211120 173816 211126 173828
rect 220081 173825 220093 173828
rect 220127 173825 220139 173859
rect 243262 173856 243268 173868
rect 220081 173819 220139 173825
rect 221660 173828 243268 173856
rect 219342 173748 219348 173800
rect 219400 173788 219406 173800
rect 221660 173788 221688 173828
rect 243262 173816 243268 173828
rect 243320 173816 243326 173868
rect 246298 173816 246304 173868
rect 246356 173856 246362 173868
rect 253842 173856 253848 173868
rect 246356 173828 253848 173856
rect 246356 173816 246362 173828
rect 253842 173816 253848 173828
rect 253900 173816 253906 173868
rect 320450 173816 320456 173868
rect 320508 173856 320514 173868
rect 409874 173856 409880 173868
rect 320508 173828 409880 173856
rect 320508 173816 320514 173828
rect 409874 173816 409880 173828
rect 409932 173816 409938 173868
rect 219400 173760 221688 173788
rect 221737 173791 221795 173797
rect 219400 173748 219406 173760
rect 221737 173757 221749 173791
rect 221783 173788 221795 173791
rect 241882 173788 241888 173800
rect 221783 173760 241888 173788
rect 221783 173757 221795 173760
rect 221737 173751 221795 173757
rect 241882 173748 241888 173760
rect 241940 173748 241946 173800
rect 246942 173748 246948 173800
rect 247000 173788 247006 173800
rect 254302 173788 254308 173800
rect 247000 173760 254308 173788
rect 247000 173748 247006 173760
rect 254302 173748 254308 173760
rect 254360 173748 254366 173800
rect 323302 173748 323308 173800
rect 323360 173788 323366 173800
rect 416774 173788 416780 173800
rect 323360 173760 416780 173788
rect 323360 173748 323366 173760
rect 416774 173748 416780 173760
rect 416832 173748 416838 173800
rect 122742 173680 122748 173732
rect 122800 173720 122806 173732
rect 204070 173720 204076 173732
rect 122800 173692 204076 173720
rect 122800 173680 122806 173692
rect 204070 173680 204076 173692
rect 204128 173680 204134 173732
rect 213822 173680 213828 173732
rect 213880 173720 213886 173732
rect 240870 173720 240876 173732
rect 213880 173692 240876 173720
rect 213880 173680 213886 173692
rect 240870 173680 240876 173692
rect 240928 173680 240934 173732
rect 245562 173680 245568 173732
rect 245620 173720 245626 173732
rect 253382 173720 253388 173732
rect 245620 173692 253388 173720
rect 245620 173680 245626 173692
rect 253382 173680 253388 173692
rect 253440 173680 253446 173732
rect 326154 173680 326160 173732
rect 326212 173720 326218 173732
rect 425054 173720 425060 173732
rect 326212 173692 425060 173720
rect 326212 173680 326218 173692
rect 425054 173680 425060 173692
rect 425112 173680 425118 173732
rect 118602 173612 118608 173664
rect 118660 173652 118666 173664
rect 202598 173652 202604 173664
rect 118660 173624 202604 173652
rect 118660 173612 118666 173624
rect 202598 173612 202604 173624
rect 202656 173612 202662 173664
rect 220081 173655 220139 173661
rect 220081 173621 220093 173655
rect 220127 173652 220139 173655
rect 239950 173652 239956 173664
rect 220127 173624 239956 173652
rect 220127 173621 220139 173624
rect 220081 173615 220139 173621
rect 239950 173612 239956 173624
rect 240008 173612 240014 173664
rect 242802 173612 242808 173664
rect 242860 173652 242866 173664
rect 252370 173652 252376 173664
rect 242860 173624 252376 173652
rect 242860 173612 242866 173624
rect 252370 173612 252376 173624
rect 252428 173612 252434 173664
rect 329006 173612 329012 173664
rect 329064 173652 329070 173664
rect 431954 173652 431960 173664
rect 329064 173624 431960 173652
rect 329064 173612 329070 173624
rect 431954 173612 431960 173624
rect 432012 173612 432018 173664
rect 111702 173544 111708 173596
rect 111760 173584 111766 173596
rect 199746 173584 199752 173596
rect 111760 173556 199752 173584
rect 111760 173544 111766 173556
rect 199746 173544 199752 173556
rect 199804 173544 199810 173596
rect 206922 173544 206928 173596
rect 206980 173584 206986 173596
rect 229465 173587 229523 173593
rect 229465 173584 229477 173587
rect 206980 173556 229477 173584
rect 206980 173544 206986 173556
rect 229465 173553 229477 173556
rect 229511 173553 229523 173587
rect 229465 173547 229523 173553
rect 229741 173587 229799 173593
rect 229741 173553 229753 173587
rect 229787 173584 229799 173587
rect 235166 173584 235172 173596
rect 229787 173556 235172 173584
rect 229787 173553 229799 173556
rect 229741 173547 229799 173553
rect 235166 173544 235172 173556
rect 235224 173544 235230 173596
rect 244918 173544 244924 173596
rect 244976 173584 244982 173596
rect 252922 173584 252928 173596
rect 244976 173556 252928 173584
rect 244976 173544 244982 173556
rect 252922 173544 252928 173556
rect 252980 173544 252986 173596
rect 331950 173544 331956 173596
rect 332008 173584 332014 173596
rect 438854 173584 438860 173596
rect 332008 173556 438860 173584
rect 332008 173544 332014 173556
rect 438854 173544 438860 173556
rect 438912 173544 438918 173596
rect 35158 173476 35164 173528
rect 35216 173516 35222 173528
rect 168098 173516 168104 173528
rect 35216 173488 168104 173516
rect 35216 173476 35222 173488
rect 168098 173476 168104 173488
rect 168156 173476 168162 173528
rect 204162 173476 204168 173528
rect 204220 173516 204226 173528
rect 229649 173519 229707 173525
rect 229649 173516 229661 173519
rect 204220 173488 229661 173516
rect 204220 173476 204226 173488
rect 229649 173485 229661 173488
rect 229695 173485 229707 173519
rect 229649 173479 229707 173485
rect 241422 173476 241428 173528
rect 241480 173516 241486 173528
rect 251910 173516 251916 173528
rect 241480 173488 251916 173516
rect 241480 173476 241486 173488
rect 251910 173476 251916 173488
rect 251968 173476 251974 173528
rect 299477 173519 299535 173525
rect 299477 173485 299489 173519
rect 299523 173516 299535 173519
rect 309045 173519 309103 173525
rect 309045 173516 309057 173519
rect 299523 173488 309057 173516
rect 299523 173485 299535 173488
rect 299477 173479 299535 173485
rect 309045 173485 309057 173488
rect 309091 173485 309103 173519
rect 309045 173479 309103 173485
rect 334802 173476 334808 173528
rect 334860 173516 334866 173528
rect 445754 173516 445760 173528
rect 334860 173488 445760 173516
rect 334860 173476 334866 173488
rect 445754 173476 445760 173488
rect 445812 173476 445818 173528
rect 29638 173408 29644 173460
rect 29696 173448 29702 173460
rect 165246 173448 165252 173460
rect 29696 173420 165252 173448
rect 29696 173408 29702 173420
rect 165246 173408 165252 173420
rect 165304 173408 165310 173460
rect 201402 173408 201408 173460
rect 201460 173448 201466 173460
rect 201460 173420 229692 173448
rect 201460 173408 201466 173420
rect 19978 173340 19984 173392
rect 20036 173380 20042 173392
rect 161382 173380 161388 173392
rect 20036 173352 161388 173380
rect 20036 173340 20042 173352
rect 161382 173340 161388 173352
rect 161440 173340 161446 173392
rect 202782 173340 202788 173392
rect 202840 173380 202846 173392
rect 229557 173383 229615 173389
rect 229557 173380 229569 173383
rect 202840 173352 229569 173380
rect 202840 173340 202846 173352
rect 229557 173349 229569 173352
rect 229603 173349 229615 173383
rect 229664 173380 229692 173420
rect 235258 173408 235264 173460
rect 235316 173448 235322 173460
rect 248046 173448 248052 173460
rect 235316 173420 248052 173448
rect 235316 173408 235322 173420
rect 248046 173408 248052 173420
rect 248104 173408 248110 173460
rect 248322 173408 248328 173460
rect 248380 173448 248386 173460
rect 254762 173448 254768 173460
rect 248380 173420 254768 173448
rect 248380 173408 248386 173420
rect 254762 173408 254768 173420
rect 254820 173408 254826 173460
rect 337654 173408 337660 173460
rect 337712 173448 337718 173460
rect 452654 173448 452660 173460
rect 337712 173420 452660 173448
rect 337712 173408 337718 173420
rect 452654 173408 452660 173420
rect 452712 173408 452718 173460
rect 235626 173380 235632 173392
rect 229664 173352 235632 173380
rect 229557 173343 229615 173349
rect 235626 173340 235632 173352
rect 235684 173340 235690 173392
rect 238662 173340 238668 173392
rect 238720 173380 238726 173392
rect 250990 173380 250996 173392
rect 238720 173352 250996 173380
rect 238720 173340 238726 173352
rect 250990 173340 250996 173352
rect 251048 173340 251054 173392
rect 309045 173383 309103 173389
rect 309045 173349 309057 173383
rect 309091 173380 309103 173383
rect 312538 173380 312544 173392
rect 309091 173352 312544 173380
rect 309091 173349 309103 173352
rect 309045 173343 309103 173349
rect 312538 173340 312544 173352
rect 312596 173340 312602 173392
rect 316696 173352 321784 173380
rect 28258 173272 28264 173324
rect 28316 173312 28322 173324
rect 164786 173312 164792 173324
rect 28316 173284 164792 173312
rect 28316 173272 28322 173284
rect 164786 173272 164792 173284
rect 164844 173272 164850 173324
rect 200022 173272 200028 173324
rect 200080 173312 200086 173324
rect 229741 173315 229799 173321
rect 229741 173312 229753 173315
rect 200080 173284 229753 173312
rect 200080 173272 200086 173284
rect 229741 173281 229753 173284
rect 229787 173281 229799 173315
rect 229741 173275 229799 173281
rect 229833 173315 229891 173321
rect 229833 173281 229845 173315
rect 229879 173312 229891 173315
rect 234525 173315 234583 173321
rect 234525 173312 234537 173315
rect 229879 173284 234537 173312
rect 229879 173281 229891 173284
rect 229833 173275 229891 173281
rect 234525 173281 234537 173284
rect 234571 173281 234583 173315
rect 234525 173275 234583 173281
rect 235902 173272 235908 173324
rect 235960 173312 235966 173324
rect 249518 173312 249524 173324
rect 235960 173284 249524 173312
rect 235960 173272 235966 173284
rect 249518 173272 249524 173284
rect 249576 173272 249582 173324
rect 273438 173272 273444 173324
rect 273496 173312 273502 173324
rect 287698 173312 287704 173324
rect 273496 173284 287704 173312
rect 273496 173272 273502 173284
rect 287698 173272 287704 173284
rect 287756 173272 287762 173324
rect 299477 173315 299535 173321
rect 299477 173312 299489 173315
rect 287808 173284 299489 173312
rect 18598 173204 18604 173256
rect 18656 173244 18662 173256
rect 160922 173244 160928 173256
rect 18656 173216 160928 173244
rect 18656 173204 18662 173216
rect 160922 173204 160928 173216
rect 160980 173204 160986 173256
rect 197262 173204 197268 173256
rect 197320 173244 197326 173256
rect 229373 173247 229431 173253
rect 229373 173244 229385 173247
rect 197320 173216 229385 173244
rect 197320 173204 197326 173216
rect 229373 173213 229385 173216
rect 229419 173213 229431 173247
rect 229373 173207 229431 173213
rect 229649 173247 229707 173253
rect 229649 173213 229661 173247
rect 229695 173244 229707 173247
rect 237098 173244 237104 173256
rect 229695 173216 237104 173244
rect 229695 173213 229707 173216
rect 229649 173207 229707 173213
rect 237098 173204 237104 173216
rect 237156 173204 237162 173256
rect 237282 173204 237288 173256
rect 237340 173244 237346 173256
rect 250530 173244 250536 173256
rect 237340 173216 250536 173244
rect 237340 173204 237346 173216
rect 250530 173204 250536 173216
rect 250588 173204 250594 173256
rect 262490 173204 262496 173256
rect 262548 173244 262554 173256
rect 266538 173244 266544 173256
rect 262548 173216 266544 173244
rect 262548 173204 262554 173216
rect 266538 173204 266544 173216
rect 266596 173204 266602 173256
rect 281166 173204 281172 173256
rect 281224 173244 281230 173256
rect 287808 173244 287836 173284
rect 299477 173281 299489 173284
rect 299523 173281 299535 173315
rect 299477 173275 299535 173281
rect 281224 173216 287836 173244
rect 281224 173204 281230 173216
rect 288342 173204 288348 173256
rect 288400 173244 288406 173256
rect 288400 173216 299520 173244
rect 288400 173204 288406 173216
rect 10318 173136 10324 173188
rect 10376 173176 10382 173188
rect 157610 173176 157616 173188
rect 10376 173148 157616 173176
rect 10376 173136 10382 173148
rect 157610 173136 157616 173148
rect 157668 173136 157674 173188
rect 194410 173136 194416 173188
rect 194468 173176 194474 173188
rect 232774 173176 232780 173188
rect 194468 173148 232780 173176
rect 194468 173136 194474 173148
rect 232774 173136 232780 173148
rect 232832 173136 232838 173188
rect 239309 173179 239367 173185
rect 239309 173145 239321 173179
rect 239355 173176 239367 173179
rect 249058 173176 249064 173188
rect 239355 173148 249064 173176
rect 239355 173145 239367 173148
rect 239309 173139 239367 173145
rect 249058 173136 249064 173148
rect 249116 173136 249122 173188
rect 251082 173136 251088 173188
rect 251140 173176 251146 173188
rect 255774 173176 255780 173188
rect 251140 173148 255780 173176
rect 251140 173136 251146 173148
rect 255774 173136 255780 173148
rect 255832 173136 255838 173188
rect 263870 173136 263876 173188
rect 263928 173176 263934 173188
rect 266998 173176 267004 173188
rect 263928 173148 267004 173176
rect 263928 173136 263934 173148
rect 266998 173136 267004 173148
rect 267056 173136 267062 173188
rect 299492 173185 299520 173216
rect 299477 173179 299535 173185
rect 299477 173145 299489 173179
rect 299523 173145 299535 173179
rect 299477 173139 299535 173145
rect 304261 173179 304319 173185
rect 304261 173145 304273 173179
rect 304307 173176 304319 173179
rect 316696 173176 316724 173352
rect 317506 173204 317512 173256
rect 317564 173244 317570 173256
rect 317564 173216 321600 173244
rect 317564 173204 317570 173216
rect 304307 173148 316724 173176
rect 304307 173145 304319 173148
rect 304261 173139 304319 173145
rect 217870 173068 217876 173120
rect 217928 173108 217934 173120
rect 242342 173108 242348 173120
rect 217928 173080 242348 173108
rect 217928 173068 217934 173080
rect 242342 173068 242348 173080
rect 242400 173068 242406 173120
rect 261938 173068 261944 173120
rect 261996 173108 262002 173120
rect 265250 173108 265256 173120
rect 261996 173080 265256 173108
rect 261996 173068 262002 173080
rect 265250 173068 265256 173080
rect 265308 173068 265314 173120
rect 267734 173068 267740 173120
rect 267792 173108 267798 173120
rect 268930 173108 268936 173120
rect 267792 173080 268936 173108
rect 267792 173068 267798 173080
rect 268930 173068 268936 173080
rect 268988 173068 268994 173120
rect 274910 173068 274916 173120
rect 274968 173108 274974 173120
rect 275830 173108 275836 173120
rect 274968 173080 275836 173108
rect 274968 173068 274974 173080
rect 275830 173068 275836 173080
rect 275888 173068 275894 173120
rect 277762 173068 277768 173120
rect 277820 173108 277826 173120
rect 278682 173108 278688 173120
rect 277820 173080 278688 173108
rect 277820 173068 277826 173080
rect 278682 173068 278688 173080
rect 278740 173068 278746 173120
rect 280706 173068 280712 173120
rect 280764 173108 280770 173120
rect 281350 173108 281356 173120
rect 280764 173080 281356 173108
rect 280764 173068 280770 173080
rect 281350 173068 281356 173080
rect 281408 173068 281414 173120
rect 281626 173068 281632 173120
rect 281684 173108 281690 173120
rect 282822 173108 282828 173120
rect 281684 173080 282828 173108
rect 281684 173068 281690 173080
rect 282822 173068 282828 173080
rect 282880 173068 282886 173120
rect 321572 173108 321600 173216
rect 321756 173176 321784 173352
rect 340506 173340 340512 173392
rect 340564 173380 340570 173392
rect 459554 173380 459560 173392
rect 340564 173352 459560 173380
rect 340564 173340 340570 173352
rect 459554 173340 459560 173352
rect 459612 173340 459618 173392
rect 331306 173312 331312 173324
rect 327552 173284 331312 173312
rect 324682 173204 324688 173256
rect 324740 173244 324746 173256
rect 325602 173244 325608 173256
rect 324740 173216 325608 173244
rect 324740 173204 324746 173216
rect 325602 173204 325608 173216
rect 325660 173204 325666 173256
rect 325694 173204 325700 173256
rect 325752 173244 325758 173256
rect 326890 173244 326896 173256
rect 325752 173216 326896 173244
rect 325752 173204 325758 173216
rect 326890 173204 326896 173216
rect 326948 173204 326954 173256
rect 327552 173176 327580 173284
rect 331306 173272 331312 173284
rect 331364 173272 331370 173324
rect 343450 173272 343456 173324
rect 343508 173312 343514 173324
rect 467834 173312 467840 173324
rect 343508 173284 467840 173312
rect 343508 173272 343514 173284
rect 467834 173272 467840 173284
rect 467892 173272 467898 173324
rect 330478 173204 330484 173256
rect 330536 173244 330542 173256
rect 331122 173244 331128 173256
rect 330536 173216 331128 173244
rect 330536 173204 330542 173216
rect 331122 173204 331128 173216
rect 331180 173204 331186 173256
rect 333330 173204 333336 173256
rect 333388 173244 333394 173256
rect 333882 173244 333888 173256
rect 333388 173216 333888 173244
rect 333388 173204 333394 173216
rect 333882 173204 333888 173216
rect 333940 173204 333946 173256
rect 337194 173204 337200 173256
rect 337252 173244 337258 173256
rect 337930 173244 337936 173256
rect 337252 173216 337936 173244
rect 337252 173204 337258 173216
rect 337930 173204 337936 173216
rect 337988 173204 337994 173256
rect 338574 173204 338580 173256
rect 338632 173244 338638 173256
rect 339218 173244 339224 173256
rect 338632 173216 339224 173244
rect 338632 173204 338638 173216
rect 339218 173204 339224 173216
rect 339276 173204 339282 173256
rect 340046 173204 340052 173256
rect 340104 173244 340110 173256
rect 340690 173244 340696 173256
rect 340104 173216 340696 173244
rect 340104 173204 340110 173216
rect 340690 173204 340696 173216
rect 340748 173204 340754 173256
rect 349154 173204 349160 173256
rect 349212 173244 349218 173256
rect 354585 173247 354643 173253
rect 349212 173216 354536 173244
rect 349212 173204 349218 173216
rect 321756 173148 327580 173176
rect 327626 173136 327632 173188
rect 327684 173176 327690 173188
rect 328362 173176 328368 173188
rect 327684 173148 328368 173176
rect 327684 173136 327690 173148
rect 328362 173136 328368 173148
rect 328420 173136 328426 173188
rect 328546 173136 328552 173188
rect 328604 173176 328610 173188
rect 329650 173176 329656 173188
rect 328604 173148 329656 173176
rect 328604 173136 328610 173148
rect 329650 173136 329656 173148
rect 329708 173136 329714 173188
rect 330018 173136 330024 173188
rect 330076 173176 330082 173188
rect 330938 173176 330944 173188
rect 330076 173148 330944 173176
rect 330076 173136 330082 173148
rect 330938 173136 330944 173148
rect 330996 173136 331002 173188
rect 331398 173136 331404 173188
rect 331456 173176 331462 173188
rect 332410 173176 332416 173188
rect 331456 173148 332416 173176
rect 331456 173136 331462 173148
rect 332410 173136 332416 173148
rect 332468 173136 332474 173188
rect 332870 173136 332876 173188
rect 332928 173176 332934 173188
rect 333698 173176 333704 173188
rect 332928 173148 333704 173176
rect 332928 173136 332934 173148
rect 333698 173136 333704 173148
rect 333756 173136 333762 173188
rect 335722 173136 335728 173188
rect 335780 173176 335786 173188
rect 336550 173176 336556 173188
rect 335780 173148 336556 173176
rect 335780 173136 335786 173148
rect 336550 173136 336556 173148
rect 336608 173136 336614 173188
rect 336734 173136 336740 173188
rect 336792 173176 336798 173188
rect 338022 173176 338028 173188
rect 336792 173148 338028 173176
rect 336792 173136 336798 173148
rect 338022 173136 338028 173148
rect 338080 173136 338086 173188
rect 338114 173136 338120 173188
rect 338172 173176 338178 173188
rect 339310 173176 339316 173188
rect 338172 173148 339316 173176
rect 338172 173136 338178 173148
rect 339310 173136 339316 173148
rect 339368 173136 339374 173188
rect 339586 173136 339592 173188
rect 339644 173176 339650 173188
rect 340782 173176 340788 173188
rect 339644 173148 340788 173176
rect 339644 173136 339650 173148
rect 340782 173136 340788 173148
rect 340840 173136 340846 173188
rect 342438 173136 342444 173188
rect 342496 173176 342502 173188
rect 343542 173176 343548 173188
rect 342496 173148 343548 173176
rect 342496 173136 342502 173148
rect 343542 173136 343548 173148
rect 343600 173136 343606 173188
rect 343910 173136 343916 173188
rect 343968 173176 343974 173188
rect 344830 173176 344836 173188
rect 343968 173148 344836 173176
rect 343968 173136 343974 173148
rect 344830 173136 344836 173148
rect 344888 173136 344894 173188
rect 345290 173136 345296 173188
rect 345348 173176 345354 173188
rect 346302 173176 346308 173188
rect 345348 173148 346308 173176
rect 345348 173136 345354 173148
rect 346302 173136 346308 173148
rect 346360 173136 346366 173188
rect 346762 173136 346768 173188
rect 346820 173176 346826 173188
rect 347590 173176 347596 173188
rect 346820 173148 347596 173176
rect 346820 173136 346826 173148
rect 347590 173136 347596 173148
rect 347648 173136 347654 173188
rect 348234 173136 348240 173188
rect 348292 173176 348298 173188
rect 349062 173176 349068 173188
rect 348292 173148 349068 173176
rect 348292 173136 348298 173148
rect 349062 173136 349068 173148
rect 349120 173136 349126 173188
rect 350626 173136 350632 173188
rect 350684 173176 350690 173188
rect 351730 173176 351736 173188
rect 350684 173148 351736 173176
rect 350684 173136 350690 173148
rect 351730 173136 351736 173148
rect 351788 173136 351794 173188
rect 352006 173136 352012 173188
rect 352064 173176 352070 173188
rect 353202 173176 353208 173188
rect 352064 173148 353208 173176
rect 352064 173136 352070 173148
rect 353202 173136 353208 173148
rect 353260 173136 353266 173188
rect 354508 173176 354536 173216
rect 354585 173213 354597 173247
rect 354631 173244 354643 173247
rect 474734 173244 474740 173256
rect 354631 173216 474740 173244
rect 354631 173213 354643 173216
rect 354585 173207 354643 173213
rect 474734 173204 474740 173216
rect 474792 173204 474798 173256
rect 481634 173176 481640 173188
rect 354508 173148 481640 173176
rect 481634 173136 481640 173148
rect 481692 173136 481698 173188
rect 519078 173136 519084 173188
rect 519136 173176 519142 173188
rect 580258 173176 580264 173188
rect 519136 173148 580264 173176
rect 519136 173136 519142 173148
rect 580258 173136 580264 173148
rect 580316 173136 580322 173188
rect 402974 173108 402980 173120
rect 321572 173080 402980 173108
rect 402974 173068 402980 173080
rect 403032 173068 403038 173120
rect 214558 173000 214564 173052
rect 214616 173040 214622 173052
rect 216490 173040 216496 173052
rect 214616 173012 216496 173040
rect 214616 173000 214622 173012
rect 216490 173000 216496 173012
rect 216548 173000 216554 173052
rect 216582 173000 216588 173052
rect 216640 173040 216646 173052
rect 221737 173043 221795 173049
rect 221737 173040 221749 173043
rect 216640 173012 221749 173040
rect 216640 173000 216646 173012
rect 221737 173009 221749 173012
rect 221783 173009 221795 173043
rect 221737 173003 221795 173009
rect 234525 173043 234583 173049
rect 234525 173009 234537 173043
rect 234571 173040 234583 173043
rect 244734 173040 244740 173052
rect 234571 173012 244740 173040
rect 234571 173009 234583 173012
rect 234525 173003 234583 173009
rect 244734 173000 244740 173012
rect 244792 173000 244798 173052
rect 249702 173000 249708 173052
rect 249760 173040 249766 173052
rect 255314 173040 255320 173052
rect 249760 173012 255320 173040
rect 249760 173000 249766 173012
rect 255314 173000 255320 173012
rect 255372 173000 255378 173052
rect 299477 173043 299535 173049
rect 299477 173009 299489 173043
rect 299523 173040 299535 173043
rect 304261 173043 304319 173049
rect 304261 173040 304273 173043
rect 299523 173012 304273 173040
rect 299523 173009 299535 173012
rect 299477 173003 299535 173009
rect 304261 173009 304273 173012
rect 304307 173009 304319 173043
rect 304261 173003 304319 173009
rect 314654 173000 314660 173052
rect 314712 173040 314718 173052
rect 396074 173040 396080 173052
rect 314712 173012 396080 173040
rect 314712 173000 314718 173012
rect 396074 173000 396080 173012
rect 396132 173000 396138 173052
rect 227622 172932 227628 172984
rect 227680 172972 227686 172984
rect 246206 172972 246212 172984
rect 227680 172944 246212 172972
rect 227680 172932 227686 172944
rect 246206 172932 246212 172944
rect 246264 172932 246270 172984
rect 270586 172932 270592 172984
rect 270644 172972 270650 172984
rect 271598 172972 271604 172984
rect 270644 172944 271604 172972
rect 270644 172932 270650 172944
rect 271598 172932 271604 172944
rect 271656 172932 271662 172984
rect 272058 172932 272064 172984
rect 272116 172972 272122 172984
rect 272978 172972 272984 172984
rect 272116 172944 272984 172972
rect 272116 172932 272122 172944
rect 272978 172932 272984 172944
rect 273036 172932 273042 172984
rect 310330 172932 310336 172984
rect 310388 172972 310394 172984
rect 385402 172972 385408 172984
rect 310388 172944 385408 172972
rect 310388 172932 310394 172944
rect 385402 172932 385408 172944
rect 385460 172932 385466 172984
rect 223482 172864 223488 172916
rect 223540 172904 223546 172916
rect 229373 172907 229431 172913
rect 223540 172876 228956 172904
rect 223540 172864 223546 172876
rect 228928 172768 228956 172876
rect 229373 172873 229385 172907
rect 229419 172904 229431 172907
rect 234246 172904 234252 172916
rect 229419 172876 234252 172904
rect 229419 172873 229431 172876
rect 229373 172867 229431 172873
rect 234246 172864 234252 172876
rect 234304 172864 234310 172916
rect 234522 172864 234528 172916
rect 234580 172904 234586 172916
rect 239309 172907 239367 172913
rect 239309 172904 239321 172907
rect 234580 172876 239321 172904
rect 234580 172864 234586 172876
rect 239309 172873 239321 172876
rect 239355 172873 239367 172907
rect 239309 172867 239367 172873
rect 239401 172907 239459 172913
rect 239401 172873 239413 172907
rect 239447 172904 239459 172907
rect 247586 172904 247592 172916
rect 239447 172876 247592 172904
rect 239447 172873 239459 172876
rect 239401 172867 239459 172873
rect 247586 172864 247592 172876
rect 247644 172864 247650 172916
rect 279234 172864 279240 172916
rect 279292 172904 279298 172916
rect 279970 172904 279976 172916
rect 279292 172876 279976 172904
rect 279292 172864 279298 172876
rect 279970 172864 279976 172876
rect 280028 172864 280034 172916
rect 307478 172864 307484 172916
rect 307536 172904 307542 172916
rect 307536 172876 374040 172904
rect 307536 172864 307542 172876
rect 229002 172796 229008 172848
rect 229060 172836 229066 172848
rect 246666 172836 246672 172848
rect 229060 172808 246672 172836
rect 229060 172796 229066 172808
rect 246666 172796 246672 172808
rect 246724 172796 246730 172848
rect 346394 172796 346400 172848
rect 346452 172836 346458 172848
rect 354585 172839 354643 172845
rect 354585 172836 354597 172839
rect 346452 172808 354597 172836
rect 346452 172796 346458 172808
rect 354585 172805 354597 172808
rect 354631 172805 354643 172839
rect 354585 172799 354643 172805
rect 354858 172796 354864 172848
rect 354916 172836 354922 172848
rect 355962 172836 355968 172848
rect 354916 172808 355968 172836
rect 354916 172796 354922 172808
rect 355962 172796 355968 172808
rect 356020 172796 356026 172848
rect 356330 172796 356336 172848
rect 356388 172836 356394 172848
rect 357342 172836 357348 172848
rect 356388 172808 357348 172836
rect 356388 172796 356394 172808
rect 357342 172796 357348 172808
rect 357400 172796 357406 172848
rect 357802 172796 357808 172848
rect 357860 172836 357866 172848
rect 358722 172836 358728 172848
rect 357860 172808 358728 172836
rect 357860 172796 357866 172808
rect 358722 172796 358728 172808
rect 358780 172796 358786 172848
rect 359182 172796 359188 172848
rect 359240 172836 359246 172848
rect 360102 172836 360108 172848
rect 359240 172808 360108 172836
rect 359240 172796 359246 172808
rect 360102 172796 360108 172808
rect 360160 172796 360166 172848
rect 360654 172796 360660 172848
rect 360712 172836 360718 172848
rect 361482 172836 361488 172848
rect 360712 172808 361488 172836
rect 360712 172796 360718 172808
rect 361482 172796 361488 172808
rect 361540 172796 361546 172848
rect 361574 172796 361580 172848
rect 361632 172836 361638 172848
rect 362770 172836 362776 172848
rect 361632 172808 362776 172836
rect 361632 172796 361638 172808
rect 362770 172796 362776 172808
rect 362828 172796 362834 172848
rect 363046 172796 363052 172848
rect 363104 172836 363110 172848
rect 364058 172836 364064 172848
rect 363104 172808 364064 172836
rect 363104 172796 363110 172808
rect 364058 172796 364064 172808
rect 364116 172796 364122 172848
rect 364518 172796 364524 172848
rect 364576 172836 364582 172848
rect 365438 172836 365444 172848
rect 364576 172808 365444 172836
rect 364576 172796 364582 172808
rect 365438 172796 365444 172808
rect 365496 172796 365502 172848
rect 365898 172796 365904 172848
rect 365956 172836 365962 172848
rect 366910 172836 366916 172848
rect 365956 172808 366916 172836
rect 365956 172796 365962 172808
rect 366910 172796 366916 172808
rect 366968 172796 366974 172848
rect 367370 172796 367376 172848
rect 367428 172836 367434 172848
rect 368290 172836 368296 172848
rect 367428 172808 368296 172836
rect 367428 172796 367434 172808
rect 368290 172796 368296 172808
rect 368348 172796 368354 172848
rect 368750 172796 368756 172848
rect 368808 172836 368814 172848
rect 369670 172836 369676 172848
rect 368808 172808 369676 172836
rect 368808 172796 368814 172808
rect 369670 172796 369676 172808
rect 369728 172796 369734 172848
rect 370222 172796 370228 172848
rect 370280 172836 370286 172848
rect 371050 172836 371056 172848
rect 370280 172808 371056 172836
rect 370280 172796 370286 172808
rect 371050 172796 371056 172808
rect 371108 172796 371114 172848
rect 371694 172796 371700 172848
rect 371752 172836 371758 172848
rect 372522 172836 372528 172848
rect 371752 172808 372528 172836
rect 371752 172796 371758 172808
rect 372522 172796 372528 172808
rect 372580 172796 372586 172848
rect 372614 172796 372620 172848
rect 372672 172836 372678 172848
rect 373902 172836 373908 172848
rect 372672 172808 373908 172836
rect 372672 172796 372678 172808
rect 373902 172796 373908 172808
rect 373960 172796 373966 172848
rect 229833 172771 229891 172777
rect 229833 172768 229845 172771
rect 228928 172740 229845 172768
rect 229833 172737 229845 172740
rect 229879 172737 229891 172771
rect 229833 172731 229891 172737
rect 232498 172728 232504 172780
rect 232556 172768 232562 172780
rect 245194 172768 245200 172780
rect 232556 172740 245200 172768
rect 232556 172728 232562 172740
rect 245194 172728 245200 172740
rect 245252 172728 245258 172780
rect 256602 172728 256608 172780
rect 256660 172768 256666 172780
rect 258166 172768 258172 172780
rect 256660 172740 258172 172768
rect 256660 172728 256666 172740
rect 258166 172728 258172 172740
rect 258224 172728 258230 172780
rect 265342 172728 265348 172780
rect 265400 172768 265406 172780
rect 266170 172768 266176 172780
rect 265400 172740 266176 172768
rect 265400 172728 265406 172740
rect 266170 172728 266176 172740
rect 266228 172728 266234 172780
rect 266814 172728 266820 172780
rect 266872 172768 266878 172780
rect 267642 172768 267648 172780
rect 266872 172740 267648 172768
rect 266872 172728 266878 172740
rect 267642 172728 267648 172740
rect 267700 172728 267706 172780
rect 268194 172728 268200 172780
rect 268252 172768 268258 172780
rect 269022 172768 269028 172780
rect 268252 172740 269028 172768
rect 268252 172728 268258 172740
rect 269022 172728 269028 172740
rect 269080 172728 269086 172780
rect 269206 172728 269212 172780
rect 269264 172768 269270 172780
rect 270218 172768 270224 172780
rect 269264 172740 270224 172768
rect 269264 172728 269270 172740
rect 270218 172728 270224 172740
rect 270276 172728 270282 172780
rect 276382 172728 276388 172780
rect 276440 172768 276446 172780
rect 277118 172768 277124 172780
rect 276440 172740 277124 172768
rect 276440 172728 276446 172740
rect 277118 172728 277124 172740
rect 277176 172728 277182 172780
rect 321830 172728 321836 172780
rect 321888 172768 321894 172780
rect 322842 172768 322848 172780
rect 321888 172740 322848 172768
rect 321888 172728 321894 172740
rect 322842 172728 322848 172740
rect 322900 172728 322906 172780
rect 340966 172728 340972 172780
rect 341024 172768 341030 172780
rect 342070 172768 342076 172780
rect 341024 172740 342076 172768
rect 341024 172728 341030 172740
rect 342070 172728 342076 172740
rect 342128 172728 342134 172780
rect 353478 172728 353484 172780
rect 353536 172768 353542 172780
rect 354490 172768 354496 172780
rect 353536 172740 354496 172768
rect 353536 172728 353542 172740
rect 354490 172728 354496 172740
rect 354548 172728 354554 172780
rect 354766 172728 354772 172780
rect 354824 172768 354830 172780
rect 355410 172768 355416 172780
rect 354824 172740 355416 172768
rect 354824 172728 354830 172740
rect 355410 172728 355416 172740
rect 355468 172728 355474 172780
rect 360194 172728 360200 172780
rect 360252 172768 360258 172780
rect 361390 172768 361396 172780
rect 360252 172740 361396 172768
rect 360252 172728 360258 172740
rect 361390 172728 361396 172740
rect 361448 172728 361454 172780
rect 373074 172728 373080 172780
rect 373132 172768 373138 172780
rect 373810 172768 373816 172780
rect 373132 172740 373816 172768
rect 373132 172728 373138 172740
rect 373810 172728 373816 172740
rect 373868 172728 373874 172780
rect 374012 172768 374040 172876
rect 374086 172864 374092 172916
rect 374144 172904 374150 172916
rect 375190 172904 375196 172916
rect 374144 172876 375196 172904
rect 374144 172864 374150 172876
rect 375190 172864 375196 172876
rect 375248 172864 375254 172916
rect 375466 172864 375472 172916
rect 375524 172904 375530 172916
rect 376570 172904 376576 172916
rect 375524 172876 376576 172904
rect 375524 172864 375530 172876
rect 376570 172864 376576 172876
rect 376628 172864 376634 172916
rect 376938 172864 376944 172916
rect 376996 172904 377002 172916
rect 377950 172904 377956 172916
rect 376996 172876 377956 172904
rect 376996 172864 377002 172876
rect 377950 172864 377956 172876
rect 378008 172864 378014 172916
rect 378410 172864 378416 172916
rect 378468 172904 378474 172916
rect 379330 172904 379336 172916
rect 378468 172876 379336 172904
rect 378468 172864 378474 172876
rect 379330 172864 379336 172876
rect 379388 172864 379394 172916
rect 374546 172796 374552 172848
rect 374604 172836 374610 172848
rect 375098 172836 375104 172848
rect 374604 172808 375104 172836
rect 374604 172796 374610 172808
rect 375098 172796 375104 172808
rect 375156 172796 375162 172848
rect 378318 172768 378324 172780
rect 374012 172740 378324 172768
rect 378318 172728 378324 172740
rect 378376 172728 378382 172780
rect 231118 172660 231124 172712
rect 231176 172700 231182 172712
rect 239401 172703 239459 172709
rect 239401 172700 239413 172703
rect 231176 172672 239413 172700
rect 231176 172660 231182 172672
rect 239401 172669 239413 172672
rect 239447 172669 239459 172703
rect 239401 172663 239459 172669
rect 243078 172660 243084 172712
rect 243136 172700 243142 172712
rect 243538 172700 243544 172712
rect 243136 172672 243544 172700
rect 243136 172660 243142 172672
rect 243538 172660 243544 172672
rect 243596 172660 243602 172712
rect 253842 172660 253848 172712
rect 253900 172700 253906 172712
rect 256694 172700 256700 172712
rect 253900 172672 256700 172700
rect 253900 172660 253906 172672
rect 256694 172660 256700 172672
rect 256752 172660 256758 172712
rect 229557 172635 229615 172641
rect 229557 172601 229569 172635
rect 229603 172632 229615 172635
rect 236638 172632 236644 172644
rect 229603 172604 236644 172632
rect 229603 172601 229615 172604
rect 229557 172595 229615 172601
rect 236638 172592 236644 172604
rect 236696 172592 236702 172644
rect 255222 172592 255228 172644
rect 255280 172632 255286 172644
rect 257706 172632 257712 172644
rect 255280 172604 257712 172632
rect 255280 172592 255286 172604
rect 257706 172592 257712 172604
rect 257764 172592 257770 172644
rect 261478 172592 261484 172644
rect 261536 172632 261542 172644
rect 262858 172632 262864 172644
rect 261536 172604 262864 172632
rect 261536 172592 261542 172604
rect 262858 172592 262864 172604
rect 262916 172592 262922 172644
rect 262950 172592 262956 172644
rect 263008 172632 263014 172644
rect 264238 172632 264244 172644
rect 263008 172604 264244 172632
rect 263008 172592 263014 172604
rect 264238 172592 264244 172604
rect 264296 172592 264302 172644
rect 265802 172592 265808 172644
rect 265860 172632 265866 172644
rect 268378 172632 268384 172644
rect 265860 172604 268384 172632
rect 265860 172592 265866 172604
rect 268378 172592 268384 172604
rect 268436 172592 268442 172644
rect 275370 172592 275376 172644
rect 275428 172632 275434 172644
rect 278038 172632 278044 172644
rect 275428 172604 278044 172632
rect 275428 172592 275434 172604
rect 278038 172592 278044 172604
rect 278096 172592 278102 172644
rect 278774 172592 278780 172644
rect 278832 172632 278838 172644
rect 280062 172632 280068 172644
rect 278832 172604 280068 172632
rect 278832 172592 278838 172604
rect 280062 172592 280068 172604
rect 280120 172592 280126 172644
rect 280154 172592 280160 172644
rect 280212 172632 280218 172644
rect 281442 172632 281448 172644
rect 280212 172604 281448 172632
rect 280212 172592 280218 172604
rect 281442 172592 281448 172604
rect 281500 172592 281506 172644
rect 283558 172592 283564 172644
rect 283616 172632 283622 172644
rect 290458 172632 290464 172644
rect 283616 172604 290464 172632
rect 283616 172592 283622 172604
rect 290458 172592 290464 172604
rect 290516 172592 290522 172644
rect 291194 172592 291200 172644
rect 291252 172632 291258 172644
rect 292390 172632 292396 172644
rect 291252 172604 292396 172632
rect 291252 172592 291258 172604
rect 292390 172592 292396 172604
rect 292448 172592 292454 172644
rect 292666 172592 292672 172644
rect 292724 172632 292730 172644
rect 293770 172632 293776 172644
rect 292724 172604 293776 172632
rect 292724 172592 292730 172604
rect 293770 172592 293776 172604
rect 293828 172592 293834 172644
rect 294506 172592 294512 172644
rect 294564 172632 294570 172644
rect 295242 172632 295248 172644
rect 294564 172604 295248 172632
rect 294564 172592 294570 172604
rect 295242 172592 295248 172604
rect 295300 172592 295306 172644
rect 295518 172592 295524 172644
rect 295576 172632 295582 172644
rect 296530 172632 296536 172644
rect 295576 172604 296536 172632
rect 295576 172592 295582 172604
rect 296530 172592 296536 172604
rect 296588 172592 296594 172644
rect 296990 172592 296996 172644
rect 297048 172632 297054 172644
rect 297910 172632 297916 172644
rect 297048 172604 297916 172632
rect 297048 172592 297054 172604
rect 297910 172592 297916 172604
rect 297968 172592 297974 172644
rect 298830 172592 298836 172644
rect 298888 172632 298894 172644
rect 299382 172632 299388 172644
rect 298888 172604 299388 172632
rect 298888 172592 298894 172604
rect 299382 172592 299388 172604
rect 299440 172592 299446 172644
rect 299842 172592 299848 172644
rect 299900 172632 299906 172644
rect 300578 172632 300584 172644
rect 299900 172604 300584 172632
rect 299900 172592 299906 172604
rect 300578 172592 300584 172604
rect 300636 172592 300642 172644
rect 302694 172592 302700 172644
rect 302752 172632 302758 172644
rect 303338 172632 303344 172644
rect 302752 172604 303344 172632
rect 302752 172592 302758 172604
rect 303338 172592 303344 172604
rect 303396 172592 303402 172644
rect 305546 172592 305552 172644
rect 305604 172632 305610 172644
rect 306098 172632 306104 172644
rect 305604 172604 306104 172632
rect 305604 172592 305610 172604
rect 306098 172592 306104 172604
rect 306156 172592 306162 172644
rect 307018 172592 307024 172644
rect 307076 172632 307082 172644
rect 307570 172632 307576 172644
rect 307076 172604 307576 172632
rect 307076 172592 307082 172604
rect 307570 172592 307576 172604
rect 307628 172592 307634 172644
rect 327074 172592 327080 172644
rect 327132 172632 327138 172644
rect 328178 172632 328184 172644
rect 327132 172604 328184 172632
rect 327132 172592 327138 172604
rect 328178 172592 328184 172604
rect 328236 172592 328242 172644
rect 334342 172592 334348 172644
rect 334400 172632 334406 172644
rect 335170 172632 335176 172644
rect 334400 172604 335176 172632
rect 334400 172592 334406 172604
rect 335170 172592 335176 172604
rect 335228 172592 335234 172644
rect 383654 172592 383660 172644
rect 383712 172632 383718 172644
rect 384942 172632 384948 172644
rect 383712 172604 384948 172632
rect 383712 172592 383718 172604
rect 384942 172592 384948 172604
rect 385000 172592 385006 172644
rect 385034 172592 385040 172644
rect 385092 172632 385098 172644
rect 386322 172632 386328 172644
rect 385092 172604 386328 172632
rect 385092 172592 385098 172604
rect 386322 172592 386328 172604
rect 386380 172592 386386 172644
rect 386506 172592 386512 172644
rect 386564 172632 386570 172644
rect 387702 172632 387708 172644
rect 386564 172604 387708 172632
rect 386564 172592 386570 172604
rect 387702 172592 387708 172604
rect 387760 172592 387766 172644
rect 387978 172592 387984 172644
rect 388036 172632 388042 172644
rect 389082 172632 389088 172644
rect 388036 172604 389088 172632
rect 388036 172592 388042 172604
rect 389082 172592 389088 172604
rect 389140 172592 389146 172644
rect 389358 172592 389364 172644
rect 389416 172632 389422 172644
rect 390462 172632 390468 172644
rect 389416 172604 390468 172632
rect 389416 172592 389422 172604
rect 390462 172592 390468 172604
rect 390520 172592 390526 172644
rect 215938 172524 215944 172576
rect 215996 172564 216002 172576
rect 217962 172564 217968 172576
rect 215996 172536 217968 172564
rect 215996 172524 216002 172536
rect 217962 172524 217968 172536
rect 218020 172524 218026 172576
rect 229465 172567 229523 172573
rect 229465 172533 229477 172567
rect 229511 172564 229523 172567
rect 238018 172564 238024 172576
rect 229511 172536 238024 172564
rect 229511 172533 229523 172536
rect 229465 172527 229523 172533
rect 238018 172524 238024 172536
rect 238076 172524 238082 172576
rect 243538 172524 243544 172576
rect 243596 172564 243602 172576
rect 248598 172564 248604 172576
rect 243596 172536 248604 172564
rect 243596 172524 243602 172536
rect 248598 172524 248604 172536
rect 248656 172524 248662 172576
rect 254578 172524 254584 172576
rect 254636 172564 254642 172576
rect 256234 172564 256240 172576
rect 254636 172536 256240 172564
rect 254636 172524 254642 172536
rect 256234 172524 256240 172536
rect 256292 172524 256298 172576
rect 260098 172524 260104 172576
rect 260156 172564 260162 172576
rect 260926 172564 260932 172576
rect 260156 172536 260932 172564
rect 260156 172524 260162 172536
rect 260926 172524 260932 172536
rect 260984 172524 260990 172576
rect 261018 172524 261024 172576
rect 261076 172564 261082 172576
rect 262122 172564 262128 172576
rect 261076 172536 262128 172564
rect 261076 172524 261082 172536
rect 262122 172524 262128 172536
rect 262180 172524 262186 172576
rect 283098 172524 283104 172576
rect 283156 172564 283162 172576
rect 284202 172564 284208 172576
rect 283156 172536 284208 172564
rect 283156 172524 283162 172536
rect 284202 172524 284208 172536
rect 284260 172524 284266 172576
rect 284478 172524 284484 172576
rect 284536 172564 284542 172576
rect 285490 172564 285496 172576
rect 284536 172536 285496 172564
rect 284536 172524 284542 172536
rect 285490 172524 285496 172536
rect 285548 172524 285554 172576
rect 285950 172524 285956 172576
rect 286008 172564 286014 172576
rect 286962 172564 286968 172576
rect 286008 172536 286968 172564
rect 286008 172524 286014 172536
rect 286962 172524 286968 172536
rect 287020 172524 287026 172576
rect 287330 172524 287336 172576
rect 287388 172564 287394 172576
rect 288342 172564 288348 172576
rect 287388 172536 288348 172564
rect 287388 172524 287394 172536
rect 288342 172524 288348 172536
rect 288400 172524 288406 172576
rect 288802 172524 288808 172576
rect 288860 172564 288866 172576
rect 289722 172564 289728 172576
rect 288860 172536 289728 172564
rect 288860 172524 288866 172536
rect 289722 172524 289728 172536
rect 289780 172524 289786 172576
rect 290274 172524 290280 172576
rect 290332 172564 290338 172576
rect 291102 172564 291108 172576
rect 290332 172536 291108 172564
rect 290332 172524 290338 172536
rect 291102 172524 291108 172536
rect 291160 172524 291166 172576
rect 291654 172524 291660 172576
rect 291712 172564 291718 172576
rect 292482 172564 292488 172576
rect 291712 172536 292488 172564
rect 291712 172524 291718 172536
rect 292482 172524 292488 172536
rect 292540 172524 292546 172576
rect 293126 172524 293132 172576
rect 293184 172564 293190 172576
rect 293862 172564 293868 172576
rect 293184 172536 293868 172564
rect 293184 172524 293190 172536
rect 293862 172524 293868 172536
rect 293920 172524 293926 172576
rect 294046 172524 294052 172576
rect 294104 172564 294110 172576
rect 295058 172564 295064 172576
rect 294104 172536 295064 172564
rect 294104 172524 294110 172536
rect 295058 172524 295064 172536
rect 295116 172524 295122 172576
rect 295978 172524 295984 172576
rect 296036 172564 296042 172576
rect 296622 172564 296628 172576
rect 296036 172536 296628 172564
rect 296036 172524 296042 172536
rect 296622 172524 296628 172536
rect 296680 172524 296686 172576
rect 297450 172524 297456 172576
rect 297508 172564 297514 172576
rect 298002 172564 298008 172576
rect 297508 172536 298008 172564
rect 297508 172524 297514 172536
rect 298002 172524 298008 172536
rect 298060 172524 298066 172576
rect 298370 172524 298376 172576
rect 298428 172564 298434 172576
rect 299198 172564 299204 172576
rect 298428 172536 299204 172564
rect 298428 172524 298434 172536
rect 299198 172524 299204 172536
rect 299256 172524 299262 172576
rect 300302 172524 300308 172576
rect 300360 172564 300366 172576
rect 300762 172564 300768 172576
rect 300360 172536 300768 172564
rect 300360 172524 300366 172536
rect 300762 172524 300768 172536
rect 300820 172524 300826 172576
rect 301222 172524 301228 172576
rect 301280 172564 301286 172576
rect 302050 172564 302056 172576
rect 301280 172536 302056 172564
rect 301280 172524 301286 172536
rect 302050 172524 302056 172536
rect 302108 172524 302114 172576
rect 302234 172524 302240 172576
rect 302292 172564 302298 172576
rect 303430 172564 303436 172576
rect 302292 172536 303436 172564
rect 302292 172524 302298 172536
rect 303430 172524 303436 172536
rect 303488 172524 303494 172576
rect 303614 172524 303620 172576
rect 303672 172564 303678 172576
rect 304810 172564 304816 172576
rect 303672 172536 304816 172564
rect 303672 172524 303678 172536
rect 304810 172524 304816 172536
rect 304868 172524 304874 172576
rect 305086 172524 305092 172576
rect 305144 172564 305150 172576
rect 306190 172564 306196 172576
rect 305144 172536 306196 172564
rect 305144 172524 305150 172536
rect 306190 172524 306196 172536
rect 306248 172524 306254 172576
rect 306558 172524 306564 172576
rect 306616 172564 306622 172576
rect 307662 172564 307668 172576
rect 306616 172536 307668 172564
rect 306616 172524 306622 172536
rect 307662 172524 307668 172536
rect 307720 172524 307726 172576
rect 307938 172524 307944 172576
rect 307996 172564 308002 172576
rect 308950 172564 308956 172576
rect 307996 172536 308956 172564
rect 307996 172524 308002 172536
rect 308950 172524 308956 172536
rect 309008 172524 309014 172576
rect 309410 172524 309416 172576
rect 309468 172564 309474 172576
rect 310422 172564 310428 172576
rect 309468 172536 310428 172564
rect 309468 172524 309474 172536
rect 310422 172524 310428 172536
rect 310480 172524 310486 172576
rect 310790 172524 310796 172576
rect 310848 172564 310854 172576
rect 311710 172564 311716 172576
rect 310848 172536 311716 172564
rect 310848 172524 310854 172536
rect 311710 172524 311716 172536
rect 311768 172524 311774 172576
rect 313274 172524 313280 172576
rect 313332 172564 313338 172576
rect 314562 172564 314568 172576
rect 313332 172536 314568 172564
rect 313332 172524 313338 172536
rect 314562 172524 314568 172536
rect 314620 172524 314626 172576
rect 315114 172524 315120 172576
rect 315172 172564 315178 172576
rect 315850 172564 315856 172576
rect 315172 172536 315856 172564
rect 315172 172524 315178 172536
rect 315850 172524 315856 172536
rect 315908 172524 315914 172576
rect 316126 172524 316132 172576
rect 316184 172564 316190 172576
rect 317322 172564 317328 172576
rect 316184 172536 317328 172564
rect 316184 172524 316190 172536
rect 317322 172524 317328 172536
rect 317380 172524 317386 172576
rect 318978 172524 318984 172576
rect 319036 172564 319042 172576
rect 320082 172564 320088 172576
rect 319036 172536 320088 172564
rect 319036 172524 319042 172536
rect 320082 172524 320088 172536
rect 320140 172524 320146 172576
rect 379790 172524 379796 172576
rect 379848 172564 379854 172576
rect 380710 172564 380716 172576
rect 379848 172536 380716 172564
rect 379848 172524 379854 172536
rect 380710 172524 380716 172536
rect 380768 172524 380774 172576
rect 381262 172524 381268 172576
rect 381320 172564 381326 172576
rect 382090 172564 382096 172576
rect 381320 172536 382096 172564
rect 381320 172524 381326 172536
rect 382090 172524 382096 172536
rect 382148 172524 382154 172576
rect 382642 172524 382648 172576
rect 382700 172564 382706 172576
rect 383562 172564 383568 172576
rect 382700 172536 383568 172564
rect 382700 172524 382706 172536
rect 383562 172524 383568 172536
rect 383620 172524 383626 172576
rect 384114 172524 384120 172576
rect 384172 172564 384178 172576
rect 384850 172564 384856 172576
rect 384172 172536 384856 172564
rect 384172 172524 384178 172536
rect 384850 172524 384856 172536
rect 384908 172524 384914 172576
rect 385586 172524 385592 172576
rect 385644 172564 385650 172576
rect 386230 172564 386236 172576
rect 385644 172536 386236 172564
rect 385644 172524 385650 172536
rect 386230 172524 386236 172536
rect 386288 172524 386294 172576
rect 386966 172524 386972 172576
rect 387024 172564 387030 172576
rect 387610 172564 387616 172576
rect 387024 172536 387616 172564
rect 387024 172524 387030 172536
rect 387610 172524 387616 172536
rect 387668 172524 387674 172576
rect 388438 172524 388444 172576
rect 388496 172564 388502 172576
rect 388990 172564 388996 172576
rect 388496 172536 388996 172564
rect 388496 172524 388502 172536
rect 388990 172524 388996 172536
rect 389048 172524 389054 172576
rect 163498 172496 163504 172508
rect 163459 172468 163504 172496
rect 163498 172456 163504 172468
rect 163556 172456 163562 172508
rect 185118 172456 185124 172508
rect 185176 172496 185182 172508
rect 185394 172496 185400 172508
rect 185176 172468 185400 172496
rect 185176 172456 185182 172468
rect 185394 172456 185400 172468
rect 185452 172456 185458 172508
rect 223853 172499 223911 172505
rect 223853 172465 223865 172499
rect 223899 172496 223911 172499
rect 224218 172496 224224 172508
rect 223899 172468 224224 172496
rect 223899 172465 223911 172468
rect 223853 172459 223911 172465
rect 224218 172456 224224 172468
rect 224276 172456 224282 172508
rect 126882 171844 126888 171896
rect 126940 171884 126946 171896
rect 205910 171884 205916 171896
rect 126940 171856 205916 171884
rect 126940 171844 126946 171856
rect 205910 171844 205916 171856
rect 205968 171844 205974 171896
rect 114462 171776 114468 171828
rect 114520 171816 114526 171828
rect 200666 171816 200672 171828
rect 114520 171788 200672 171816
rect 114520 171776 114526 171788
rect 200666 171776 200672 171788
rect 200724 171776 200730 171828
rect 349614 171776 349620 171828
rect 349672 171816 349678 171828
rect 483014 171816 483020 171828
rect 349672 171788 483020 171816
rect 349672 171776 349678 171788
rect 483014 171776 483020 171788
rect 483072 171776 483078 171828
rect 225506 171096 225512 171148
rect 225564 171136 225570 171148
rect 226058 171136 226064 171148
rect 225564 171108 226064 171136
rect 225564 171096 225570 171108
rect 226058 171096 226064 171108
rect 226116 171096 226122 171148
rect 154574 171028 154580 171080
rect 154632 171068 154638 171080
rect 155310 171068 155316 171080
rect 154632 171040 155316 171068
rect 154632 171028 154638 171040
rect 155310 171028 155316 171040
rect 155368 171028 155374 171080
rect 169754 171028 169760 171080
rect 169812 171068 169818 171080
rect 170582 171068 170588 171080
rect 169812 171040 170588 171068
rect 169812 171028 169818 171040
rect 170582 171028 170588 171040
rect 170640 171028 170646 171080
rect 171134 171028 171140 171080
rect 171192 171068 171198 171080
rect 172054 171068 172060 171080
rect 171192 171040 172060 171068
rect 171192 171028 171198 171040
rect 172054 171028 172060 171040
rect 172112 171028 172118 171080
rect 175366 171028 175372 171080
rect 175424 171068 175430 171080
rect 175918 171068 175924 171080
rect 175424 171040 175924 171068
rect 175424 171028 175430 171040
rect 175918 171028 175924 171040
rect 175976 171028 175982 171080
rect 176654 171028 176660 171080
rect 176712 171068 176718 171080
rect 177114 171068 177120 171080
rect 176712 171040 177120 171068
rect 176712 171028 176718 171040
rect 177114 171028 177120 171040
rect 177172 171028 177178 171080
rect 178034 171028 178040 171080
rect 178092 171068 178098 171080
rect 178310 171068 178316 171080
rect 178092 171040 178316 171068
rect 178092 171028 178098 171040
rect 178310 171028 178316 171040
rect 178368 171028 178374 171080
rect 179414 171028 179420 171080
rect 179472 171068 179478 171080
rect 179874 171068 179880 171080
rect 179472 171040 179880 171068
rect 179472 171028 179478 171040
rect 179874 171028 179880 171040
rect 179932 171028 179938 171080
rect 186406 171028 186412 171080
rect 186464 171068 186470 171080
rect 186958 171068 186964 171080
rect 186464 171040 186964 171068
rect 186464 171028 186470 171040
rect 186958 171028 186964 171040
rect 187016 171028 187022 171080
rect 187786 171028 187792 171080
rect 187844 171068 187850 171080
rect 188430 171068 188436 171080
rect 187844 171040 188436 171068
rect 187844 171028 187850 171040
rect 188430 171028 188436 171040
rect 188488 171028 188494 171080
rect 189074 171028 189080 171080
rect 189132 171068 189138 171080
rect 189350 171068 189356 171080
rect 189132 171040 189356 171068
rect 189132 171028 189138 171040
rect 189350 171028 189356 171040
rect 189408 171028 189414 171080
rect 190546 171028 190552 171080
rect 190604 171068 190610 171080
rect 191190 171068 191196 171080
rect 190604 171040 191196 171068
rect 190604 171028 190610 171040
rect 191190 171028 191196 171040
rect 191248 171028 191254 171080
rect 191926 171028 191932 171080
rect 191984 171068 191990 171080
rect 192662 171068 192668 171080
rect 191984 171040 192668 171068
rect 191984 171028 191990 171040
rect 192662 171028 192668 171040
rect 192720 171028 192726 171080
rect 193306 171028 193312 171080
rect 193364 171068 193370 171080
rect 194134 171068 194140 171080
rect 193364 171040 194140 171068
rect 193364 171028 193370 171040
rect 194134 171028 194140 171040
rect 194192 171028 194198 171080
rect 194686 171028 194692 171080
rect 194744 171068 194750 171080
rect 195606 171068 195612 171080
rect 194744 171040 195612 171068
rect 194744 171028 194750 171040
rect 195606 171028 195612 171040
rect 195664 171028 195670 171080
rect 202966 171028 202972 171080
rect 203024 171068 203030 171080
rect 203150 171068 203156 171080
rect 203024 171040 203156 171068
rect 203024 171028 203030 171040
rect 203150 171028 203156 171040
rect 203208 171028 203214 171080
rect 204254 171028 204260 171080
rect 204312 171068 204318 171080
rect 205174 171068 205180 171080
rect 204312 171040 205180 171068
rect 204312 171028 204318 171040
rect 205174 171028 205180 171040
rect 205232 171028 205238 171080
rect 208394 171028 208400 171080
rect 208452 171068 208458 171080
rect 209038 171068 209044 171080
rect 208452 171040 209044 171068
rect 208452 171028 208458 171040
rect 209038 171028 209044 171040
rect 209096 171028 209102 171080
rect 211246 171028 211252 171080
rect 211304 171068 211310 171080
rect 211798 171068 211804 171080
rect 211304 171040 211804 171068
rect 211304 171028 211310 171040
rect 211798 171028 211804 171040
rect 211856 171028 211862 171080
rect 214006 171028 214012 171080
rect 214064 171068 214070 171080
rect 214742 171068 214748 171080
rect 214064 171040 214748 171068
rect 214064 171028 214070 171040
rect 214742 171028 214748 171040
rect 214800 171028 214806 171080
rect 227806 171028 227812 171080
rect 227864 171068 227870 171080
rect 228542 171068 228548 171080
rect 227864 171040 228548 171068
rect 227864 171028 227870 171040
rect 228542 171028 228548 171040
rect 228600 171028 228606 171080
rect 229186 171028 229192 171080
rect 229244 171068 229250 171080
rect 230014 171068 230020 171080
rect 229244 171040 230020 171068
rect 229244 171028 229250 171040
rect 230014 171028 230020 171040
rect 230072 171028 230078 171080
rect 230474 171028 230480 171080
rect 230532 171068 230538 171080
rect 230934 171068 230940 171080
rect 230532 171040 230940 171068
rect 230532 171028 230538 171040
rect 230934 171028 230940 171040
rect 230992 171028 230998 171080
rect 237466 171028 237472 171080
rect 237524 171068 237530 171080
rect 238110 171068 238116 171080
rect 237524 171040 238116 171068
rect 237524 171028 237530 171040
rect 238110 171028 238116 171040
rect 238168 171028 238174 171080
rect 240502 171028 240508 171080
rect 240560 171068 240566 171080
rect 241146 171068 241152 171080
rect 240560 171040 241152 171068
rect 240560 171028 240566 171040
rect 241146 171028 241152 171040
rect 241204 171028 241210 171080
rect 393222 171028 393228 171080
rect 393280 171068 393286 171080
rect 579890 171068 579896 171080
rect 393280 171040 579896 171068
rect 393280 171028 393286 171040
rect 579890 171028 579896 171040
rect 579948 171028 579954 171080
rect 175274 170960 175280 171012
rect 175332 171000 175338 171012
rect 175550 171000 175556 171012
rect 175332 170972 175556 171000
rect 175332 170960 175338 170972
rect 175550 170960 175556 170972
rect 175608 170960 175614 171012
rect 176746 170960 176752 171012
rect 176804 171000 176810 171012
rect 177390 171000 177396 171012
rect 176804 170972 177396 171000
rect 176804 170960 176810 170972
rect 177390 170960 177396 170972
rect 177448 170960 177454 171012
rect 179506 170960 179512 171012
rect 179564 171000 179570 171012
rect 180150 171000 180156 171012
rect 179564 170972 180156 171000
rect 179564 170960 179570 170972
rect 180150 170960 180156 170972
rect 180208 170960 180214 171012
rect 186314 170960 186320 171012
rect 186372 171000 186378 171012
rect 186590 171000 186596 171012
rect 186372 170972 186596 171000
rect 186372 170960 186378 170972
rect 186590 170960 186596 170972
rect 186648 170960 186654 171012
rect 189166 170960 189172 171012
rect 189224 171000 189230 171012
rect 189902 171000 189908 171012
rect 189224 170972 189908 171000
rect 189224 170960 189230 170972
rect 189902 170960 189908 170972
rect 189960 170960 189966 171012
rect 230566 170960 230572 171012
rect 230624 171000 230630 171012
rect 231486 171000 231492 171012
rect 230624 170972 231492 171000
rect 230624 170960 230630 170972
rect 231486 170960 231492 170972
rect 231544 170960 231550 171012
rect 218054 170484 218060 170536
rect 218112 170524 218118 170536
rect 218606 170524 218612 170536
rect 218112 170496 218612 170524
rect 218112 170484 218118 170496
rect 218606 170484 218612 170496
rect 218664 170484 218670 170536
rect 131022 170416 131028 170468
rect 131080 170456 131086 170468
rect 207014 170456 207020 170468
rect 131080 170428 207020 170456
rect 131080 170416 131086 170428
rect 207014 170416 207020 170428
rect 207072 170416 207078 170468
rect 36538 170348 36544 170400
rect 36596 170388 36602 170400
rect 169018 170388 169024 170400
rect 36596 170360 169024 170388
rect 36596 170348 36602 170360
rect 169018 170348 169024 170360
rect 169076 170348 169082 170400
rect 312262 170348 312268 170400
rect 312320 170388 312326 170400
rect 390554 170388 390560 170400
rect 312320 170360 390560 170388
rect 312320 170348 312326 170360
rect 390554 170348 390560 170360
rect 390612 170348 390618 170400
rect 187694 169396 187700 169448
rect 187752 169436 187758 169448
rect 188154 169436 188160 169448
rect 187752 169408 188160 169436
rect 187752 169396 187758 169408
rect 188154 169396 188160 169408
rect 188212 169396 188218 169448
rect 188065 169303 188123 169309
rect 188065 169269 188077 169303
rect 188111 169300 188123 169303
rect 188154 169300 188160 169312
rect 188111 169272 188160 169300
rect 188111 169269 188123 169272
rect 188065 169263 188123 169269
rect 188154 169260 188160 169272
rect 188212 169260 188218 169312
rect 159082 169124 159088 169176
rect 159140 169164 159146 169176
rect 159266 169164 159272 169176
rect 159140 169136 159272 169164
rect 159140 169124 159146 169136
rect 159266 169124 159272 169136
rect 159324 169124 159330 169176
rect 137922 169056 137928 169108
rect 137980 169096 137986 169108
rect 210234 169096 210240 169108
rect 137980 169068 210240 169096
rect 137980 169056 137986 169068
rect 210234 169056 210240 169068
rect 210292 169056 210298 169108
rect 217042 169056 217048 169108
rect 217100 169096 217106 169108
rect 217226 169096 217232 169108
rect 217100 169068 217232 169096
rect 217100 169056 217106 169068
rect 217226 169056 217232 169068
rect 217284 169056 217290 169108
rect 96522 168988 96528 169040
rect 96580 169028 96586 169040
rect 193490 169028 193496 169040
rect 96580 169000 193496 169028
rect 96580 168988 96586 169000
rect 193490 168988 193496 169000
rect 193548 168988 193554 169040
rect 350626 168988 350632 169040
rect 350684 169028 350690 169040
rect 485774 169028 485780 169040
rect 350684 169000 485780 169028
rect 350684 168988 350690 169000
rect 485774 168988 485780 169000
rect 485832 168988 485838 169040
rect 157426 168308 157432 168360
rect 157484 168348 157490 168360
rect 158254 168348 158260 168360
rect 157484 168320 158260 168348
rect 157484 168308 157490 168320
rect 158254 168308 158260 168320
rect 158312 168308 158318 168360
rect 158806 168308 158812 168360
rect 158864 168348 158870 168360
rect 159726 168348 159732 168360
rect 158864 168320 159732 168348
rect 158864 168308 158870 168320
rect 159726 168308 159732 168320
rect 159784 168308 159790 168360
rect 212626 167900 212632 167952
rect 212684 167940 212690 167952
rect 213270 167940 213276 167952
rect 212684 167912 213276 167940
rect 212684 167900 212690 167912
rect 213270 167900 213276 167912
rect 213328 167900 213334 167952
rect 194594 167832 194600 167884
rect 194652 167872 194658 167884
rect 195054 167872 195060 167884
rect 194652 167844 195060 167872
rect 194652 167832 194658 167844
rect 195054 167832 195060 167844
rect 195112 167832 195118 167884
rect 142062 167696 142068 167748
rect 142120 167736 142126 167748
rect 211706 167736 211712 167748
rect 142120 167708 211712 167736
rect 142120 167696 142126 167708
rect 211706 167696 211712 167708
rect 211764 167696 211770 167748
rect 32398 167628 32404 167680
rect 32456 167668 32462 167680
rect 167638 167668 167644 167680
rect 32456 167640 167644 167668
rect 32456 167628 32462 167640
rect 167638 167628 167644 167640
rect 167696 167628 167702 167680
rect 178126 167628 178132 167680
rect 178184 167668 178190 167680
rect 178862 167668 178868 167680
rect 178184 167640 178868 167668
rect 178184 167628 178190 167640
rect 178862 167628 178868 167640
rect 178920 167628 178926 167680
rect 352006 167628 352012 167680
rect 352064 167668 352070 167680
rect 489914 167668 489920 167680
rect 352064 167640 489920 167668
rect 352064 167628 352070 167640
rect 489914 167628 489920 167640
rect 489972 167628 489978 167680
rect 209866 167424 209872 167476
rect 209924 167464 209930 167476
rect 210326 167464 210332 167476
rect 209924 167436 210332 167464
rect 209924 167424 209930 167436
rect 210326 167424 210332 167436
rect 210384 167424 210390 167476
rect 207198 167356 207204 167408
rect 207256 167396 207262 167408
rect 208026 167396 208032 167408
rect 207256 167368 208032 167396
rect 207256 167356 207262 167368
rect 208026 167356 208032 167368
rect 208084 167356 208090 167408
rect 156230 167016 156236 167068
rect 156288 167056 156294 167068
rect 156874 167056 156880 167068
rect 156288 167028 156880 167056
rect 156288 167016 156294 167028
rect 156874 167016 156880 167028
rect 156932 167016 156938 167068
rect 201494 167016 201500 167068
rect 201552 167056 201558 167068
rect 201678 167056 201684 167068
rect 201552 167028 201684 167056
rect 201552 167016 201558 167028
rect 201678 167016 201684 167028
rect 201736 167016 201742 167068
rect 215294 167016 215300 167068
rect 215352 167056 215358 167068
rect 215478 167056 215484 167068
rect 215352 167028 215484 167056
rect 215352 167016 215358 167028
rect 215478 167016 215484 167028
rect 215536 167016 215542 167068
rect 256878 166948 256884 167000
rect 256936 166988 256942 167000
rect 257062 166988 257068 167000
rect 256936 166960 257068 166988
rect 256936 166948 256942 166960
rect 257062 166948 257068 166960
rect 257120 166948 257126 167000
rect 133782 166336 133788 166388
rect 133840 166376 133846 166388
rect 208486 166376 208492 166388
rect 133840 166348 208492 166376
rect 133840 166336 133846 166348
rect 208486 166336 208492 166348
rect 208544 166336 208550 166388
rect 38562 166268 38568 166320
rect 38620 166308 38626 166320
rect 169938 166308 169944 166320
rect 38620 166280 169944 166308
rect 38620 166268 38626 166280
rect 169938 166268 169944 166280
rect 169996 166268 170002 166320
rect 353386 166268 353392 166320
rect 353444 166308 353450 166320
rect 494054 166308 494060 166320
rect 353444 166280 494060 166308
rect 353444 166268 353450 166280
rect 494054 166268 494060 166280
rect 494112 166268 494118 166320
rect 3234 165520 3240 165572
rect 3292 165560 3298 165572
rect 153102 165560 153108 165572
rect 3292 165532 153108 165560
rect 3292 165520 3298 165532
rect 153102 165520 153108 165532
rect 153160 165520 153166 165572
rect 174078 165316 174084 165368
rect 174136 165356 174142 165368
rect 174538 165356 174544 165368
rect 174136 165328 174544 165356
rect 174136 165316 174142 165328
rect 174538 165316 174544 165328
rect 174596 165316 174602 165368
rect 144822 164840 144828 164892
rect 144880 164880 144886 164892
rect 212718 164880 212724 164892
rect 144880 164852 212724 164880
rect 144880 164840 144886 164852
rect 212718 164840 212724 164852
rect 212776 164840 212782 164892
rect 354766 164840 354772 164892
rect 354824 164880 354830 164892
rect 496814 164880 496820 164892
rect 354824 164852 496820 164880
rect 354824 164840 354830 164852
rect 496814 164840 496820 164852
rect 496872 164840 496878 164892
rect 181162 164228 181168 164280
rect 181220 164268 181226 164280
rect 181714 164268 181720 164280
rect 181220 164240 181720 164268
rect 181220 164228 181226 164240
rect 181714 164228 181720 164240
rect 181772 164228 181778 164280
rect 182450 164228 182456 164280
rect 182508 164268 182514 164280
rect 183186 164268 183192 164280
rect 182508 164240 183192 164268
rect 182508 164228 182514 164240
rect 183186 164228 183192 164240
rect 183244 164228 183250 164280
rect 183922 164228 183928 164280
rect 183980 164268 183986 164280
rect 184474 164268 184480 164280
rect 183980 164240 184480 164268
rect 183980 164228 183986 164240
rect 184474 164228 184480 164240
rect 184532 164228 184538 164280
rect 168374 164160 168380 164212
rect 168432 164200 168438 164212
rect 168650 164200 168656 164212
rect 168432 164172 168656 164200
rect 168432 164160 168438 164172
rect 168650 164160 168656 164172
rect 168708 164160 168714 164212
rect 172422 164160 172428 164212
rect 172480 164200 172486 164212
rect 172698 164200 172704 164212
rect 172480 164172 172704 164200
rect 172480 164160 172486 164172
rect 172698 164160 172704 164172
rect 172756 164160 172762 164212
rect 206002 164200 206008 164212
rect 205963 164172 206008 164200
rect 206002 164160 206008 164172
rect 206060 164160 206066 164212
rect 216950 164160 216956 164212
rect 217008 164200 217014 164212
rect 217042 164200 217048 164212
rect 217008 164172 217048 164200
rect 217008 164160 217014 164172
rect 217042 164160 217048 164172
rect 217100 164160 217106 164212
rect 240502 164200 240508 164212
rect 240463 164172 240508 164200
rect 240502 164160 240508 164172
rect 240560 164160 240566 164212
rect 256786 164160 256792 164212
rect 256844 164200 256850 164212
rect 257062 164200 257068 164212
rect 256844 164172 257068 164200
rect 256844 164160 256850 164172
rect 257062 164160 257068 164172
rect 257120 164160 257126 164212
rect 385218 164200 385224 164212
rect 385179 164172 385224 164200
rect 385218 164160 385224 164172
rect 385276 164160 385282 164212
rect 148962 163548 148968 163600
rect 149020 163588 149026 163600
rect 214098 163588 214104 163600
rect 149020 163560 214104 163588
rect 149020 163548 149026 163560
rect 214098 163548 214104 163560
rect 214156 163548 214162 163600
rect 31018 163480 31024 163532
rect 31076 163520 31082 163532
rect 165798 163520 165804 163532
rect 31076 163492 165804 163520
rect 31076 163480 31082 163492
rect 165798 163480 165804 163492
rect 165856 163480 165862 163532
rect 357158 163480 357164 163532
rect 357216 163520 357222 163532
rect 500954 163520 500960 163532
rect 357216 163492 500960 163520
rect 357216 163480 357222 163492
rect 500954 163480 500960 163492
rect 501012 163480 501018 163532
rect 163038 162868 163044 162920
rect 163096 162908 163102 162920
rect 163501 162911 163559 162917
rect 163501 162908 163513 162911
rect 163096 162880 163513 162908
rect 163096 162868 163102 162880
rect 163501 162877 163513 162880
rect 163547 162877 163559 162911
rect 223850 162908 223856 162920
rect 223811 162880 223856 162908
rect 163501 162871 163559 162877
rect 223850 162868 223856 162880
rect 223908 162868 223914 162920
rect 163130 162800 163136 162852
rect 163188 162840 163194 162852
rect 163314 162840 163320 162852
rect 163188 162812 163320 162840
rect 163188 162800 163194 162812
rect 163314 162800 163320 162812
rect 163372 162800 163378 162852
rect 174078 162800 174084 162852
rect 174136 162840 174142 162852
rect 174262 162840 174268 162852
rect 174136 162812 174268 162840
rect 174136 162800 174142 162812
rect 174262 162800 174268 162812
rect 174320 162800 174326 162852
rect 181162 162840 181168 162852
rect 181123 162812 181168 162840
rect 181162 162800 181168 162812
rect 181220 162800 181226 162852
rect 151722 162188 151728 162240
rect 151780 162228 151786 162240
rect 215386 162228 215392 162240
rect 151780 162200 215392 162228
rect 151780 162188 151786 162200
rect 215386 162188 215392 162200
rect 215444 162188 215450 162240
rect 21358 162120 21364 162172
rect 21416 162160 21422 162172
rect 161566 162160 161572 162172
rect 21416 162132 161572 162160
rect 21416 162120 21422 162132
rect 161566 162120 161572 162132
rect 161624 162120 161630 162172
rect 201678 162120 201684 162172
rect 201736 162120 201742 162172
rect 358538 162120 358544 162172
rect 358596 162160 358602 162172
rect 503714 162160 503720 162172
rect 358596 162132 503720 162160
rect 358596 162120 358602 162132
rect 503714 162120 503720 162132
rect 503772 162120 503778 162172
rect 201696 161968 201724 162120
rect 201678 161916 201684 161968
rect 201736 161916 201742 161968
rect 163041 161415 163099 161421
rect 163041 161381 163053 161415
rect 163087 161412 163099 161415
rect 163314 161412 163320 161424
rect 163087 161384 163320 161412
rect 163087 161381 163099 161384
rect 163041 161375 163099 161381
rect 163314 161372 163320 161384
rect 163372 161372 163378 161424
rect 225325 161415 225383 161421
rect 225325 161381 225337 161415
rect 225371 161412 225383 161415
rect 225414 161412 225420 161424
rect 225371 161384 225420 161412
rect 225371 161381 225383 161384
rect 225325 161375 225383 161381
rect 225414 161372 225420 161384
rect 225472 161372 225478 161424
rect 132402 160760 132408 160812
rect 132460 160800 132466 160812
rect 207106 160800 207112 160812
rect 132460 160772 207112 160800
rect 132460 160760 132466 160772
rect 207106 160760 207112 160772
rect 207164 160760 207170 160812
rect 55122 160692 55128 160744
rect 55180 160732 55186 160744
rect 176838 160732 176844 160744
rect 55180 160704 176844 160732
rect 55180 160692 55186 160704
rect 176838 160692 176844 160704
rect 176896 160692 176902 160744
rect 360010 160692 360016 160744
rect 360068 160732 360074 160744
rect 507854 160732 507860 160744
rect 360068 160704 507860 160732
rect 360068 160692 360074 160704
rect 507854 160692 507860 160704
rect 507912 160692 507918 160744
rect 201494 159400 201500 159452
rect 201552 159440 201558 159452
rect 201862 159440 201868 159452
rect 201552 159412 201868 159440
rect 201552 159400 201558 159412
rect 201862 159400 201868 159412
rect 201920 159400 201926 159452
rect 128262 159332 128268 159384
rect 128320 159372 128326 159384
rect 205726 159372 205732 159384
rect 128320 159344 205732 159372
rect 128320 159332 128326 159344
rect 205726 159332 205732 159344
rect 205784 159332 205790 159384
rect 361298 159332 361304 159384
rect 361356 159372 361362 159384
rect 511994 159372 512000 159384
rect 361356 159344 512000 159372
rect 361356 159332 361362 159344
rect 511994 159332 512000 159344
rect 512052 159332 512058 159384
rect 393130 158652 393136 158704
rect 393188 158692 393194 158704
rect 580166 158692 580172 158704
rect 393188 158664 580172 158692
rect 393188 158652 393194 158664
rect 580166 158652 580172 158664
rect 580224 158652 580230 158704
rect 146202 158040 146208 158092
rect 146260 158080 146266 158092
rect 212626 158080 212632 158092
rect 146260 158052 212632 158080
rect 146260 158040 146266 158052
rect 212626 158040 212632 158052
rect 212684 158040 212690 158092
rect 11698 157972 11704 158024
rect 11756 158012 11762 158024
rect 158898 158012 158904 158024
rect 11756 157984 158904 158012
rect 11756 157972 11762 157984
rect 158898 157972 158904 157984
rect 158956 157972 158962 158024
rect 198918 157496 198924 157548
rect 198976 157496 198982 157548
rect 198936 157344 198964 157496
rect 226518 157360 226524 157412
rect 226576 157400 226582 157412
rect 226702 157400 226708 157412
rect 226576 157372 226708 157400
rect 226576 157360 226582 157372
rect 226702 157360 226708 157372
rect 226760 157360 226766 157412
rect 198918 157292 198924 157344
rect 198976 157292 198982 157344
rect 385218 157332 385224 157344
rect 385179 157304 385224 157332
rect 385218 157292 385224 157304
rect 385276 157292 385282 157344
rect 139302 156680 139308 156732
rect 139360 156720 139366 156732
rect 209866 156720 209872 156732
rect 139360 156692 209872 156720
rect 139360 156680 139366 156692
rect 209866 156680 209872 156692
rect 209924 156680 209930 156732
rect 314378 156680 314384 156732
rect 314436 156720 314442 156732
rect 393314 156720 393320 156732
rect 314436 156692 393320 156720
rect 314436 156680 314442 156692
rect 393314 156680 393320 156692
rect 393372 156680 393378 156732
rect 50982 156612 50988 156664
rect 51040 156652 51046 156664
rect 175458 156652 175464 156664
rect 51040 156624 175464 156652
rect 51040 156612 51046 156624
rect 175458 156612 175464 156624
rect 175516 156612 175522 156664
rect 364058 156612 364064 156664
rect 364116 156652 364122 156664
rect 516134 156652 516140 156664
rect 364116 156624 516140 156652
rect 364116 156612 364122 156624
rect 516134 156612 516140 156624
rect 516192 156612 516198 156664
rect 240502 156312 240508 156324
rect 240463 156284 240508 156312
rect 240502 156272 240508 156284
rect 240560 156272 240566 156324
rect 150342 155252 150348 155304
rect 150400 155292 150406 155304
rect 214006 155292 214012 155304
rect 150400 155264 214012 155292
rect 150400 155252 150406 155264
rect 214006 155252 214012 155264
rect 214064 155252 214070 155304
rect 315850 155252 315856 155304
rect 315908 155292 315914 155304
rect 397454 155292 397460 155304
rect 315908 155264 397460 155292
rect 315908 155252 315914 155264
rect 397454 155252 397460 155264
rect 397512 155252 397518 155304
rect 42702 155184 42708 155236
rect 42760 155224 42766 155236
rect 171410 155224 171416 155236
rect 42760 155196 171416 155224
rect 42760 155184 42766 155196
rect 171410 155184 171416 155196
rect 171468 155184 171474 155236
rect 365438 155184 365444 155236
rect 365496 155224 365502 155236
rect 520274 155224 520280 155236
rect 365496 155196 520280 155224
rect 365496 155184 365502 155196
rect 520274 155184 520280 155196
rect 520332 155184 520338 155236
rect 206002 154612 206008 154624
rect 205963 154584 206008 154612
rect 206002 154572 206008 154584
rect 206060 154572 206066 154624
rect 210050 154572 210056 154624
rect 210108 154612 210114 154624
rect 210142 154612 210148 154624
rect 210108 154584 210148 154612
rect 210108 154572 210114 154584
rect 210142 154572 210148 154584
rect 210200 154572 210206 154624
rect 207198 154504 207204 154556
rect 207256 154544 207262 154556
rect 207474 154544 207480 154556
rect 207256 154516 207480 154544
rect 207256 154504 207262 154516
rect 207474 154504 207480 154516
rect 207532 154504 207538 154556
rect 218238 154504 218244 154556
rect 218296 154544 218302 154556
rect 218422 154544 218428 154556
rect 218296 154516 218428 154544
rect 218296 154504 218302 154516
rect 218422 154504 218428 154516
rect 218480 154504 218486 154556
rect 219526 154504 219532 154556
rect 219584 154544 219590 154556
rect 219710 154544 219716 154556
rect 219584 154516 219716 154544
rect 219584 154504 219590 154516
rect 219710 154504 219716 154516
rect 219768 154504 219774 154556
rect 256970 154504 256976 154556
rect 257028 154544 257034 154556
rect 257154 154544 257160 154556
rect 257028 154516 257160 154544
rect 257028 154504 257034 154516
rect 257154 154504 257160 154516
rect 257212 154504 257218 154556
rect 317138 153892 317144 153944
rect 317196 153932 317202 153944
rect 400306 153932 400312 153944
rect 317196 153904 400312 153932
rect 317196 153892 317202 153904
rect 400306 153892 400312 153904
rect 400364 153892 400370 153944
rect 82722 153824 82728 153876
rect 82780 153864 82786 153876
rect 188246 153864 188252 153876
rect 82780 153836 188252 153864
rect 82780 153824 82786 153836
rect 188246 153824 188252 153836
rect 188304 153824 188310 153876
rect 362678 153824 362684 153876
rect 362736 153864 362742 153876
rect 513374 153864 513380 153876
rect 362736 153836 513380 153864
rect 362736 153824 362742 153836
rect 513374 153824 513380 153836
rect 513432 153824 513438 153876
rect 183922 153348 183928 153400
rect 183980 153348 183986 153400
rect 183940 153264 183968 153348
rect 183922 153212 183928 153264
rect 183980 153212 183986 153264
rect 185210 153212 185216 153264
rect 185268 153252 185274 153264
rect 185302 153252 185308 153264
rect 185268 153224 185308 153252
rect 185268 153212 185274 153224
rect 185302 153212 185308 153224
rect 185360 153212 185366 153264
rect 318610 152532 318616 152584
rect 318668 152572 318674 152584
rect 404354 152572 404360 152584
rect 318668 152544 404360 152572
rect 318668 152532 318674 152544
rect 404354 152532 404360 152544
rect 404412 152532 404418 152584
rect 85482 152464 85488 152516
rect 85540 152504 85546 152516
rect 189258 152504 189264 152516
rect 85540 152476 189264 152504
rect 85540 152464 85546 152476
rect 189258 152464 189264 152476
rect 189316 152464 189322 152516
rect 366818 152464 366824 152516
rect 366876 152504 366882 152516
rect 524414 152504 524420 152516
rect 366876 152476 524420 152504
rect 366876 152464 366882 152476
rect 524414 152464 524420 152476
rect 524472 152464 524478 152516
rect 163038 151824 163044 151836
rect 162999 151796 163044 151824
rect 163038 151784 163044 151796
rect 163096 151784 163102 151836
rect 225322 151824 225328 151836
rect 225283 151796 225328 151824
rect 225322 151784 225328 151796
rect 225380 151784 225386 151836
rect 378134 151784 378140 151836
rect 378192 151824 378198 151836
rect 378318 151824 378324 151836
rect 378192 151796 378324 151824
rect 378192 151784 378198 151796
rect 378318 151784 378324 151796
rect 378376 151784 378382 151836
rect 223758 151756 223764 151768
rect 223719 151728 223764 151756
rect 223758 151716 223764 151728
rect 223816 151716 223822 151768
rect 319898 151104 319904 151156
rect 319956 151144 319962 151156
rect 408494 151144 408500 151156
rect 319956 151116 408500 151144
rect 319956 151104 319962 151116
rect 408494 151104 408500 151116
rect 408552 151104 408558 151156
rect 89622 151036 89628 151088
rect 89680 151076 89686 151088
rect 190638 151076 190644 151088
rect 89680 151048 190644 151076
rect 89680 151036 89686 151048
rect 190638 151036 190644 151048
rect 190696 151036 190702 151088
rect 279878 151036 279884 151088
rect 279936 151076 279942 151088
rect 309134 151076 309140 151088
rect 279936 151048 309140 151076
rect 279936 151036 279942 151048
rect 309134 151036 309140 151048
rect 309192 151036 309198 151088
rect 368198 151036 368204 151088
rect 368256 151076 368262 151088
rect 528554 151076 528560 151088
rect 368256 151048 528560 151076
rect 368256 151036 368262 151048
rect 528554 151036 528560 151048
rect 528612 151036 528618 151088
rect 321370 149744 321376 149796
rect 321428 149784 321434 149796
rect 411254 149784 411260 149796
rect 321428 149756 411260 149784
rect 321428 149744 321434 149756
rect 411254 149744 411260 149756
rect 411312 149744 411318 149796
rect 92382 149676 92388 149728
rect 92440 149716 92446 149728
rect 192018 149716 192024 149728
rect 92440 149688 192024 149716
rect 92440 149676 92446 149688
rect 192018 149676 192024 149688
rect 192076 149676 192082 149728
rect 369578 149676 369584 149728
rect 369636 149716 369642 149728
rect 531314 149716 531320 149728
rect 369636 149688 531320 149716
rect 369636 149676 369642 149688
rect 531314 149676 531320 149688
rect 531372 149676 531378 149728
rect 322658 148384 322664 148436
rect 322716 148424 322722 148436
rect 415394 148424 415400 148436
rect 322716 148396 415400 148424
rect 322716 148384 322722 148396
rect 415394 148384 415400 148396
rect 415452 148384 415458 148436
rect 99282 148316 99288 148368
rect 99340 148356 99346 148368
rect 194778 148356 194784 148368
rect 99340 148328 194784 148356
rect 99340 148316 99346 148328
rect 194778 148316 194784 148328
rect 194836 148316 194842 148368
rect 370958 148316 370964 148368
rect 371016 148356 371022 148368
rect 535454 148356 535460 148368
rect 371016 148328 535460 148356
rect 371016 148316 371022 148328
rect 535454 148316 535460 148328
rect 535512 148316 535518 148368
rect 156230 147636 156236 147688
rect 156288 147676 156294 147688
rect 156414 147676 156420 147688
rect 156288 147648 156420 147676
rect 156288 147636 156294 147648
rect 156414 147636 156420 147648
rect 156472 147636 156478 147688
rect 168558 147636 168564 147688
rect 168616 147636 168622 147688
rect 206002 147636 206008 147688
rect 206060 147636 206066 147688
rect 226518 147636 226524 147688
rect 226576 147636 226582 147688
rect 385126 147636 385132 147688
rect 385184 147676 385190 147688
rect 385310 147676 385316 147688
rect 385184 147648 385316 147676
rect 385184 147636 385190 147648
rect 385310 147636 385316 147648
rect 385368 147636 385374 147688
rect 168576 147608 168604 147636
rect 168650 147608 168656 147620
rect 168576 147580 168656 147608
rect 168650 147568 168656 147580
rect 168708 147568 168714 147620
rect 206020 147608 206048 147636
rect 206094 147608 206100 147620
rect 206020 147580 206100 147608
rect 206094 147568 206100 147580
rect 206152 147568 206158 147620
rect 226536 147608 226564 147636
rect 226610 147608 226616 147620
rect 226536 147580 226616 147608
rect 226610 147568 226616 147580
rect 226668 147568 226674 147620
rect 324130 146956 324136 147008
rect 324188 146996 324194 147008
rect 418154 146996 418160 147008
rect 324188 146968 418160 146996
rect 324188 146956 324194 146968
rect 418154 146956 418160 146968
rect 418212 146956 418218 147008
rect 103422 146888 103428 146940
rect 103480 146928 103486 146940
rect 196066 146928 196072 146940
rect 103480 146900 196072 146928
rect 103480 146888 103486 146900
rect 196066 146888 196072 146900
rect 196124 146888 196130 146940
rect 373718 146888 373724 146940
rect 373776 146928 373782 146940
rect 542354 146928 542360 146940
rect 373776 146900 542360 146928
rect 373776 146888 373782 146900
rect 542354 146888 542360 146900
rect 542412 146888 542418 146940
rect 107562 145528 107568 145580
rect 107620 145568 107626 145580
rect 197538 145568 197544 145580
rect 107620 145540 197544 145568
rect 107620 145528 107626 145540
rect 197538 145528 197544 145540
rect 197596 145528 197602 145580
rect 353110 145528 353116 145580
rect 353168 145568 353174 145580
rect 491294 145568 491300 145580
rect 353168 145540 491300 145568
rect 353168 145528 353174 145540
rect 491294 145528 491300 145540
rect 491352 145528 491358 145580
rect 181162 145024 181168 145036
rect 181123 144996 181168 145024
rect 181162 144984 181168 144996
rect 181220 144984 181226 145036
rect 193490 144848 193496 144900
rect 193548 144888 193554 144900
rect 193582 144888 193588 144900
rect 193548 144860 193588 144888
rect 193548 144848 193554 144860
rect 193582 144848 193588 144860
rect 193640 144848 193646 144900
rect 200298 144848 200304 144900
rect 200356 144888 200362 144900
rect 200390 144888 200396 144900
rect 200356 144860 200396 144888
rect 200356 144848 200362 144860
rect 200390 144848 200396 144860
rect 200448 144848 200454 144900
rect 385218 144888 385224 144900
rect 385179 144860 385224 144888
rect 385218 144848 385224 144860
rect 385276 144848 385282 144900
rect 110322 144168 110328 144220
rect 110380 144208 110386 144220
rect 194134 144208 194140 144220
rect 110380 144180 194140 144208
rect 110380 144168 110386 144180
rect 194134 144168 194140 144180
rect 194192 144168 194198 144220
rect 358630 144168 358636 144220
rect 358688 144208 358694 144220
rect 505094 144208 505100 144220
rect 358688 144180 505100 144208
rect 358688 144168 358694 144180
rect 505094 144168 505100 144180
rect 505152 144168 505158 144220
rect 158990 143528 158996 143540
rect 158951 143500 158996 143528
rect 158990 143488 158996 143500
rect 159048 143488 159054 143540
rect 163133 143531 163191 143537
rect 163133 143497 163145 143531
rect 163179 143528 163191 143531
rect 163222 143528 163228 143540
rect 163179 143500 163228 143528
rect 163179 143497 163191 143500
rect 163133 143491 163191 143497
rect 163222 143488 163228 143500
rect 163280 143488 163286 143540
rect 168374 143488 168380 143540
rect 168432 143528 168438 143540
rect 168650 143528 168656 143540
rect 168432 143500 168656 143528
rect 168432 143488 168438 143500
rect 168650 143488 168656 143500
rect 168708 143488 168714 143540
rect 179598 143528 179604 143540
rect 179559 143500 179604 143528
rect 179598 143488 179604 143500
rect 179656 143488 179662 143540
rect 181073 143531 181131 143537
rect 181073 143497 181085 143531
rect 181119 143528 181131 143531
rect 181162 143528 181168 143540
rect 181119 143500 181168 143528
rect 181119 143497 181131 143500
rect 181073 143491 181131 143497
rect 181162 143488 181168 143500
rect 181220 143488 181226 143540
rect 183833 143531 183891 143537
rect 183833 143497 183845 143531
rect 183879 143528 183891 143531
rect 183922 143528 183928 143540
rect 183879 143500 183928 143528
rect 183879 143497 183891 143500
rect 183833 143491 183891 143497
rect 183922 143488 183928 143500
rect 183980 143488 183986 143540
rect 207290 143528 207296 143540
rect 207251 143500 207296 143528
rect 207290 143488 207296 143500
rect 207348 143488 207354 143540
rect 219618 143528 219624 143540
rect 219579 143500 219624 143528
rect 219618 143488 219624 143500
rect 219676 143488 219682 143540
rect 117222 142808 117228 142860
rect 117280 142848 117286 142860
rect 201494 142848 201500 142860
rect 117280 142820 201500 142848
rect 117280 142808 117286 142820
rect 201494 142808 201500 142820
rect 201552 142808 201558 142860
rect 357250 142808 357256 142860
rect 357308 142848 357314 142860
rect 502334 142848 502340 142860
rect 357308 142820 502340 142848
rect 357308 142808 357314 142820
rect 502334 142808 502340 142820
rect 502392 142808 502398 142860
rect 223761 142171 223819 142177
rect 223761 142137 223773 142171
rect 223807 142168 223819 142171
rect 223850 142168 223856 142180
rect 223807 142140 223856 142168
rect 223807 142137 223819 142140
rect 223761 142131 223819 142137
rect 223850 142128 223856 142140
rect 223908 142128 223914 142180
rect 121362 141380 121368 141432
rect 121420 141420 121426 141432
rect 202966 141420 202972 141432
rect 121420 141392 202972 141420
rect 121420 141380 121426 141392
rect 202966 141380 202972 141392
rect 203024 141380 203030 141432
rect 355870 141380 355876 141432
rect 355928 141420 355934 141432
rect 498194 141420 498200 141432
rect 355928 141392 498200 141420
rect 355928 141380 355934 141392
rect 498194 141380 498200 141392
rect 498252 141380 498258 141432
rect 125502 140020 125508 140072
rect 125560 140060 125566 140072
rect 204530 140060 204536 140072
rect 125560 140032 204536 140060
rect 125560 140020 125566 140032
rect 204530 140020 204536 140032
rect 204588 140020 204594 140072
rect 362770 140020 362776 140072
rect 362828 140060 362834 140072
rect 512086 140060 512092 140072
rect 362828 140032 512092 140060
rect 362828 140020 362834 140032
rect 512086 140020 512092 140032
rect 512144 140020 512150 140072
rect 46842 138660 46848 138712
rect 46900 138700 46906 138712
rect 172606 138700 172612 138712
rect 46900 138672 172612 138700
rect 46900 138660 46906 138672
rect 172606 138660 172612 138672
rect 172664 138660 172670 138712
rect 361390 138660 361396 138712
rect 361448 138700 361454 138712
rect 509234 138700 509240 138712
rect 361448 138672 509240 138700
rect 361448 138660 361454 138672
rect 509234 138660 509240 138672
rect 509292 138660 509298 138712
rect 240413 138159 240471 138165
rect 240413 138125 240425 138159
rect 240459 138156 240471 138159
rect 240502 138156 240508 138168
rect 240459 138128 240508 138156
rect 240459 138125 240471 138128
rect 240413 138119 240471 138125
rect 240502 138116 240508 138128
rect 240560 138116 240566 138168
rect 157610 138048 157616 138100
rect 157668 138048 157674 138100
rect 217042 138048 217048 138100
rect 217100 138048 217106 138100
rect 243078 138088 243084 138100
rect 243004 138060 243084 138088
rect 157628 137964 157656 138048
rect 205910 137980 205916 138032
rect 205968 138020 205974 138032
rect 206094 138020 206100 138032
rect 205968 137992 206100 138020
rect 205968 137980 205974 137992
rect 206094 137980 206100 137992
rect 206152 137980 206158 138032
rect 217060 137964 217088 138048
rect 243004 138032 243032 138060
rect 243078 138048 243084 138060
rect 243136 138048 243142 138100
rect 242986 137980 242992 138032
rect 243044 137980 243050 138032
rect 256878 137980 256884 138032
rect 256936 137980 256942 138032
rect 157610 137912 157616 137964
rect 157668 137912 157674 137964
rect 217042 137912 217048 137964
rect 217100 137912 217106 137964
rect 256896 137952 256924 137980
rect 256970 137952 256976 137964
rect 256896 137924 256976 137952
rect 256970 137912 256976 137924
rect 257028 137912 257034 137964
rect 385218 137952 385224 137964
rect 385179 137924 385224 137952
rect 385218 137912 385224 137924
rect 385276 137912 385282 137964
rect 57882 137232 57888 137284
rect 57940 137272 57946 137284
rect 178218 137272 178224 137284
rect 57940 137244 178224 137272
rect 57940 137232 57946 137244
rect 178218 137232 178224 137244
rect 178276 137232 178282 137284
rect 341978 137232 341984 137284
rect 342036 137272 342042 137284
rect 462314 137272 462320 137284
rect 342036 137244 462320 137272
rect 342036 137232 342042 137244
rect 462314 137232 462320 137244
rect 462372 137232 462378 137284
rect 3326 136552 3332 136604
rect 3384 136592 3390 136604
rect 152918 136592 152924 136604
rect 3384 136564 152924 136592
rect 3384 136552 3390 136564
rect 152918 136552 152924 136564
rect 152976 136552 152982 136604
rect 344738 135872 344744 135924
rect 344796 135912 344802 135924
rect 469214 135912 469220 135924
rect 344796 135884 469220 135912
rect 344796 135872 344802 135884
rect 469214 135872 469220 135884
rect 469272 135872 469278 135924
rect 210053 135235 210111 135241
rect 210053 135201 210065 135235
rect 210099 135232 210111 135235
rect 210142 135232 210148 135244
rect 210099 135204 210148 135232
rect 210099 135201 210111 135204
rect 210053 135195 210111 135201
rect 210142 135192 210148 135204
rect 210200 135192 210206 135244
rect 256970 135192 256976 135244
rect 257028 135232 257034 135244
rect 257154 135232 257160 135244
rect 257028 135204 257160 135232
rect 257028 135192 257034 135204
rect 257154 135192 257160 135204
rect 257212 135192 257218 135244
rect 393038 135192 393044 135244
rect 393096 135232 393102 135244
rect 579890 135232 579896 135244
rect 393096 135204 579896 135232
rect 393096 135192 393102 135204
rect 579890 135192 579896 135204
rect 579948 135192 579954 135244
rect 62022 134512 62028 134564
rect 62080 134552 62086 134564
rect 179601 134555 179659 134561
rect 179601 134552 179613 134555
rect 62080 134524 179613 134552
rect 62080 134512 62086 134524
rect 179601 134521 179613 134524
rect 179647 134521 179659 134555
rect 179601 134515 179659 134521
rect 181070 134008 181076 134020
rect 181031 133980 181076 134008
rect 181070 133968 181076 133980
rect 181128 133968 181134 134020
rect 219618 134008 219624 134020
rect 219579 133980 219624 134008
rect 219618 133968 219624 133980
rect 219676 133968 219682 134020
rect 240410 133940 240416 133952
rect 240371 133912 240416 133940
rect 240410 133900 240416 133912
rect 240468 133900 240474 133952
rect 157613 133875 157671 133881
rect 157613 133841 157625 133875
rect 157659 133872 157671 133875
rect 157794 133872 157800 133884
rect 157659 133844 157800 133872
rect 157659 133841 157671 133844
rect 157613 133835 157671 133841
rect 157794 133832 157800 133844
rect 157852 133832 157858 133884
rect 181070 133872 181076 133884
rect 181031 133844 181076 133872
rect 181070 133832 181076 133844
rect 181128 133832 181134 133884
rect 219618 133832 219624 133884
rect 219676 133872 219682 133884
rect 219710 133872 219716 133884
rect 219676 133844 219716 133872
rect 219676 133832 219682 133844
rect 219710 133832 219716 133844
rect 219768 133832 219774 133884
rect 222381 133875 222439 133881
rect 222381 133841 222393 133875
rect 222427 133872 222439 133875
rect 222470 133872 222476 133884
rect 222427 133844 222476 133872
rect 222427 133841 222439 133844
rect 222381 133835 222439 133841
rect 222470 133832 222476 133844
rect 222528 133832 222534 133884
rect 343450 133152 343456 133204
rect 343508 133192 343514 133204
rect 466454 133192 466460 133204
rect 343508 133164 466460 133192
rect 343508 133152 343514 133164
rect 466454 133152 466460 133164
rect 466512 133152 466518 133204
rect 378134 132472 378140 132524
rect 378192 132512 378198 132524
rect 378318 132512 378324 132524
rect 378192 132484 378324 132512
rect 378192 132472 378198 132484
rect 378318 132472 378324 132484
rect 378376 132472 378382 132524
rect 347498 131724 347504 131776
rect 347556 131764 347562 131776
rect 477586 131764 477592 131776
rect 347556 131736 477592 131764
rect 347556 131724 347562 131736
rect 477586 131724 477592 131736
rect 477644 131724 477650 131776
rect 158993 131019 159051 131025
rect 158993 130985 159005 131019
rect 159039 131016 159051 131019
rect 159082 131016 159088 131028
rect 159039 130988 159088 131016
rect 159039 130985 159051 130988
rect 158993 130979 159051 130985
rect 159082 130976 159088 130988
rect 159140 130976 159146 131028
rect 346210 130364 346216 130416
rect 346268 130404 346274 130416
rect 473354 130404 473360 130416
rect 346268 130376 473360 130404
rect 346268 130364 346274 130376
rect 473354 130364 473360 130376
rect 473412 130364 473418 130416
rect 354490 129004 354496 129056
rect 354548 129044 354554 129056
rect 492674 129044 492680 129056
rect 354548 129016 492680 129044
rect 354548 129004 354554 129016
rect 492674 129004 492680 129016
rect 492732 129004 492738 129056
rect 156230 128324 156236 128376
rect 156288 128364 156294 128376
rect 156414 128364 156420 128376
rect 156288 128336 156420 128364
rect 156288 128324 156294 128336
rect 156414 128324 156420 128336
rect 156472 128324 156478 128376
rect 174078 128324 174084 128376
rect 174136 128364 174142 128376
rect 174262 128364 174268 128376
rect 174136 128336 174268 128364
rect 174136 128324 174142 128336
rect 174262 128324 174268 128336
rect 174320 128324 174326 128376
rect 193398 128324 193404 128376
rect 193456 128364 193462 128376
rect 193582 128364 193588 128376
rect 193456 128336 193588 128364
rect 193456 128324 193462 128336
rect 193582 128324 193588 128336
rect 193640 128324 193646 128376
rect 205726 128324 205732 128376
rect 205784 128364 205790 128376
rect 205910 128364 205916 128376
rect 205784 128336 205916 128364
rect 205784 128324 205790 128336
rect 205910 128324 205916 128336
rect 205968 128324 205974 128376
rect 239030 128324 239036 128376
rect 239088 128324 239094 128376
rect 163130 128296 163136 128308
rect 163091 128268 163136 128296
rect 163130 128256 163136 128268
rect 163188 128256 163194 128308
rect 207290 128296 207296 128308
rect 207251 128268 207296 128296
rect 207290 128256 207296 128268
rect 207348 128256 207354 128308
rect 210050 128296 210056 128308
rect 210011 128268 210056 128296
rect 210050 128256 210056 128268
rect 210108 128256 210114 128308
rect 239048 128296 239076 128324
rect 239122 128296 239128 128308
rect 239048 128268 239128 128296
rect 239122 128256 239128 128268
rect 239180 128256 239186 128308
rect 348970 127576 348976 127628
rect 349028 127616 349034 127628
rect 480254 127616 480260 127628
rect 349028 127588 480260 127616
rect 349028 127576 349034 127588
rect 480254 127576 480260 127588
rect 480312 127576 480318 127628
rect 372430 126216 372436 126268
rect 372488 126256 372494 126268
rect 538214 126256 538220 126268
rect 372488 126228 538220 126256
rect 372488 126216 372494 126228
rect 538214 126216 538220 126228
rect 538272 126216 538278 126268
rect 182358 125536 182364 125588
rect 182416 125576 182422 125588
rect 182450 125576 182456 125588
rect 182416 125548 182456 125576
rect 182416 125536 182422 125548
rect 182450 125536 182456 125548
rect 182508 125536 182514 125588
rect 196158 125576 196164 125588
rect 196119 125548 196164 125576
rect 196158 125536 196164 125548
rect 196216 125536 196222 125588
rect 197630 125576 197636 125588
rect 197591 125548 197636 125576
rect 197630 125536 197636 125548
rect 197688 125536 197694 125588
rect 216950 125536 216956 125588
rect 217008 125576 217014 125588
rect 217042 125576 217048 125588
rect 217008 125548 217048 125576
rect 217008 125536 217014 125548
rect 217042 125536 217048 125548
rect 217100 125536 217106 125588
rect 218238 125536 218244 125588
rect 218296 125576 218302 125588
rect 218422 125576 218428 125588
rect 218296 125548 218428 125576
rect 218296 125536 218302 125548
rect 218422 125536 218428 125548
rect 218480 125536 218486 125588
rect 220998 125536 221004 125588
rect 221056 125576 221062 125588
rect 221182 125576 221188 125588
rect 221056 125548 221188 125576
rect 221056 125536 221062 125548
rect 221182 125536 221188 125548
rect 221240 125536 221246 125588
rect 364150 124856 364156 124908
rect 364208 124896 364214 124908
rect 517514 124896 517520 124908
rect 364208 124868 517520 124896
rect 364208 124856 364214 124868
rect 517514 124856 517520 124868
rect 517572 124856 517578 124908
rect 183833 124287 183891 124293
rect 183833 124253 183845 124287
rect 183879 124284 183891 124287
rect 183922 124284 183928 124296
rect 183879 124256 183928 124284
rect 183879 124253 183891 124256
rect 183833 124247 183891 124253
rect 183922 124244 183928 124256
rect 183980 124244 183986 124296
rect 223761 124287 223819 124293
rect 223761 124253 223773 124287
rect 223807 124284 223819 124287
rect 223850 124284 223856 124296
rect 223807 124256 223856 124284
rect 223807 124253 223819 124256
rect 223761 124247 223819 124253
rect 223850 124244 223856 124256
rect 223908 124244 223914 124296
rect 157610 124216 157616 124228
rect 157571 124188 157616 124216
rect 157610 124176 157616 124188
rect 157668 124176 157674 124228
rect 181073 124219 181131 124225
rect 181073 124185 181085 124219
rect 181119 124216 181131 124219
rect 181162 124216 181168 124228
rect 181119 124188 181168 124216
rect 181119 124185 181131 124188
rect 181073 124179 181131 124185
rect 181162 124176 181168 124188
rect 181220 124176 181226 124228
rect 222378 124216 222384 124228
rect 222339 124188 222384 124216
rect 222378 124176 222384 124188
rect 222436 124176 222442 124228
rect 385034 124176 385040 124228
rect 385092 124216 385098 124228
rect 385310 124216 385316 124228
rect 385092 124188 385316 124216
rect 385092 124176 385098 124188
rect 385310 124176 385316 124188
rect 385368 124176 385374 124228
rect 240410 124148 240416 124160
rect 240371 124120 240416 124148
rect 240410 124108 240416 124120
rect 240468 124108 240474 124160
rect 392946 124108 392952 124160
rect 393004 124148 393010 124160
rect 579890 124148 579896 124160
rect 393004 124120 579896 124148
rect 393004 124108 393010 124120
rect 579890 124108 579896 124120
rect 579948 124108 579954 124160
rect 223758 122856 223764 122868
rect 223719 122828 223764 122856
rect 223758 122816 223764 122828
rect 223816 122816 223822 122868
rect 3326 122748 3332 122800
rect 3384 122788 3390 122800
rect 153010 122788 153016 122800
rect 3384 122760 153016 122788
rect 3384 122748 3390 122760
rect 153010 122748 153016 122760
rect 153068 122748 153074 122800
rect 158901 122791 158959 122797
rect 158901 122757 158913 122791
rect 158947 122788 158959 122791
rect 159082 122788 159088 122800
rect 158947 122760 159088 122788
rect 158947 122757 158959 122760
rect 158901 122751 158959 122757
rect 159082 122748 159088 122760
rect 159140 122748 159146 122800
rect 183830 122748 183836 122800
rect 183888 122788 183894 122800
rect 183925 122791 183983 122797
rect 183925 122788 183937 122791
rect 183888 122760 183937 122788
rect 183888 122748 183894 122760
rect 183925 122757 183937 122760
rect 183971 122757 183983 122791
rect 183925 122751 183983 122757
rect 238754 122748 238760 122800
rect 238812 122788 238818 122800
rect 239122 122788 239128 122800
rect 238812 122760 239128 122788
rect 238812 122748 238818 122760
rect 239122 122748 239128 122760
rect 239180 122748 239186 122800
rect 218333 119391 218391 119397
rect 218333 119357 218345 119391
rect 218379 119388 218391 119391
rect 218422 119388 218428 119400
rect 218379 119360 218428 119388
rect 218379 119357 218391 119360
rect 218333 119351 218391 119357
rect 218422 119348 218428 119360
rect 218480 119348 218486 119400
rect 219621 119391 219679 119397
rect 219621 119357 219633 119391
rect 219667 119388 219679 119391
rect 219710 119388 219716 119400
rect 219667 119360 219716 119388
rect 219667 119357 219679 119360
rect 219621 119351 219679 119357
rect 219710 119348 219716 119360
rect 219768 119348 219774 119400
rect 385034 119348 385040 119400
rect 385092 119388 385098 119400
rect 385092 119360 385137 119388
rect 385092 119348 385098 119360
rect 163038 118668 163044 118720
rect 163096 118708 163102 118720
rect 163222 118708 163228 118720
rect 163096 118680 163228 118708
rect 163096 118668 163102 118680
rect 163222 118668 163228 118680
rect 163280 118668 163286 118720
rect 174170 118668 174176 118720
rect 174228 118668 174234 118720
rect 205818 118668 205824 118720
rect 205876 118668 205882 118720
rect 207290 118668 207296 118720
rect 207348 118668 207354 118720
rect 226610 118668 226616 118720
rect 226668 118668 226674 118720
rect 256878 118668 256884 118720
rect 256936 118668 256942 118720
rect 174188 118640 174216 118668
rect 174262 118640 174268 118652
rect 174188 118612 174268 118640
rect 174262 118600 174268 118612
rect 174320 118600 174326 118652
rect 205836 118640 205864 118668
rect 205910 118640 205916 118652
rect 205836 118612 205916 118640
rect 205910 118600 205916 118612
rect 205968 118600 205974 118652
rect 207308 118640 207336 118668
rect 207382 118640 207388 118652
rect 207308 118612 207388 118640
rect 207382 118600 207388 118612
rect 207440 118600 207446 118652
rect 226628 118640 226656 118668
rect 226702 118640 226708 118652
rect 226628 118612 226708 118640
rect 226702 118600 226708 118612
rect 226760 118600 226766 118652
rect 256896 118640 256924 118668
rect 256970 118640 256976 118652
rect 256896 118612 256976 118640
rect 256970 118600 256976 118612
rect 257028 118600 257034 118652
rect 181162 115988 181168 116000
rect 181123 115960 181168 115988
rect 181162 115948 181168 115960
rect 181220 115948 181226 116000
rect 185118 115948 185124 116000
rect 185176 115988 185182 116000
rect 185210 115988 185216 116000
rect 185176 115960 185216 115988
rect 185176 115948 185182 115960
rect 185210 115948 185216 115960
rect 185268 115948 185274 116000
rect 196158 115988 196164 116000
rect 196119 115960 196164 115988
rect 196158 115948 196164 115960
rect 196216 115948 196222 116000
rect 197630 115988 197636 116000
rect 197591 115960 197636 115988
rect 197630 115948 197636 115960
rect 197688 115948 197694 116000
rect 223758 115948 223764 116000
rect 223816 115948 223822 116000
rect 225230 115948 225236 116000
rect 225288 115948 225294 116000
rect 163130 115920 163136 115932
rect 163091 115892 163136 115920
rect 163130 115880 163136 115892
rect 163188 115880 163194 115932
rect 222378 115880 222384 115932
rect 222436 115920 222442 115932
rect 222562 115920 222568 115932
rect 222436 115892 222568 115920
rect 222436 115880 222442 115892
rect 222562 115880 222568 115892
rect 222620 115880 222626 115932
rect 223776 115852 223804 115948
rect 223850 115852 223856 115864
rect 223776 115824 223856 115852
rect 223850 115812 223856 115824
rect 223908 115812 223914 115864
rect 225248 115852 225276 115948
rect 228082 115920 228088 115932
rect 228043 115892 228088 115920
rect 228082 115880 228088 115892
rect 228140 115880 228146 115932
rect 256970 115880 256976 115932
rect 257028 115920 257034 115932
rect 257154 115920 257160 115932
rect 257028 115892 257160 115920
rect 257028 115880 257034 115892
rect 257154 115880 257160 115892
rect 257212 115880 257218 115932
rect 225322 115852 225328 115864
rect 225248 115824 225328 115852
rect 225322 115812 225328 115824
rect 225380 115812 225386 115864
rect 168558 114520 168564 114572
rect 168616 114560 168622 114572
rect 168650 114560 168656 114572
rect 168616 114532 168656 114560
rect 168616 114520 168622 114532
rect 168650 114520 168656 114532
rect 168708 114520 168714 114572
rect 180978 114520 180984 114572
rect 181036 114560 181042 114572
rect 181165 114563 181223 114569
rect 181165 114560 181177 114563
rect 181036 114532 181177 114560
rect 181036 114520 181042 114532
rect 181165 114529 181177 114532
rect 181211 114529 181223 114563
rect 218330 114560 218336 114572
rect 218291 114532 218336 114560
rect 181165 114523 181223 114529
rect 218330 114520 218336 114532
rect 218388 114520 218394 114572
rect 219618 114560 219624 114572
rect 219579 114532 219624 114560
rect 219618 114520 219624 114532
rect 219676 114520 219682 114572
rect 240410 114560 240416 114572
rect 240371 114532 240416 114560
rect 240410 114520 240416 114532
rect 240468 114520 240474 114572
rect 185118 114492 185124 114504
rect 185079 114464 185124 114492
rect 185118 114452 185124 114464
rect 185176 114452 185182 114504
rect 180978 114424 180984 114436
rect 180939 114396 180984 114424
rect 180978 114384 180984 114396
rect 181036 114384 181042 114436
rect 158898 113200 158904 113212
rect 158859 113172 158904 113200
rect 158898 113160 158904 113172
rect 158956 113160 158962 113212
rect 183922 113160 183928 113212
rect 183980 113200 183986 113212
rect 183980 113172 184025 113200
rect 183980 113160 183986 113172
rect 378134 113160 378140 113212
rect 378192 113200 378198 113212
rect 378318 113200 378324 113212
rect 378192 113172 378324 113200
rect 378192 113160 378198 113172
rect 378318 113160 378324 113172
rect 378376 113160 378382 113212
rect 158898 113064 158904 113076
rect 158859 113036 158904 113064
rect 158898 113024 158904 113036
rect 158956 113024 158962 113076
rect 395338 111732 395344 111784
rect 395396 111772 395402 111784
rect 580166 111772 580172 111784
rect 395396 111744 580172 111772
rect 395396 111732 395402 111744
rect 580166 111732 580172 111744
rect 580224 111732 580230 111784
rect 225322 111228 225328 111240
rect 225248 111200 225328 111228
rect 225248 111172 225276 111200
rect 225322 111188 225328 111200
rect 225380 111188 225386 111240
rect 225230 111120 225236 111172
rect 225288 111120 225294 111172
rect 185121 111027 185179 111033
rect 185121 110993 185133 111027
rect 185167 111024 185179 111027
rect 185210 111024 185216 111036
rect 185167 110996 185216 111024
rect 185167 110993 185179 110996
rect 185121 110987 185179 110993
rect 185210 110984 185216 110996
rect 185268 110984 185274 111036
rect 156230 109012 156236 109064
rect 156288 109052 156294 109064
rect 156414 109052 156420 109064
rect 156288 109024 156420 109052
rect 156288 109012 156294 109024
rect 156414 109012 156420 109024
rect 156472 109012 156478 109064
rect 157610 109012 157616 109064
rect 157668 109012 157674 109064
rect 174078 109012 174084 109064
rect 174136 109052 174142 109064
rect 174262 109052 174268 109064
rect 174136 109024 174268 109052
rect 174136 109012 174142 109024
rect 174262 109012 174268 109024
rect 174320 109012 174326 109064
rect 193398 109012 193404 109064
rect 193456 109052 193462 109064
rect 193582 109052 193588 109064
rect 193456 109024 193588 109052
rect 193456 109012 193462 109024
rect 193582 109012 193588 109024
rect 193640 109012 193646 109064
rect 205726 109012 205732 109064
rect 205784 109052 205790 109064
rect 205910 109052 205916 109064
rect 205784 109024 205916 109052
rect 205784 109012 205790 109024
rect 205910 109012 205916 109024
rect 205968 109012 205974 109064
rect 157628 108984 157656 109012
rect 157702 108984 157708 108996
rect 157628 108956 157708 108984
rect 157702 108944 157708 108956
rect 157760 108944 157766 108996
rect 163130 108984 163136 108996
rect 163091 108956 163136 108984
rect 163130 108944 163136 108956
rect 163188 108944 163194 108996
rect 218330 106332 218336 106344
rect 218256 106304 218336 106332
rect 218256 106276 218284 106304
rect 218330 106292 218336 106304
rect 218388 106292 218394 106344
rect 221090 106332 221096 106344
rect 221016 106304 221096 106332
rect 221016 106276 221044 106304
rect 221090 106292 221096 106304
rect 221148 106292 221154 106344
rect 228082 106332 228088 106344
rect 228043 106304 228088 106332
rect 228082 106292 228088 106304
rect 228140 106292 228146 106344
rect 385034 106332 385040 106344
rect 384995 106304 385040 106332
rect 385034 106292 385040 106304
rect 385092 106292 385098 106344
rect 196158 106264 196164 106276
rect 196119 106236 196164 106264
rect 196158 106224 196164 106236
rect 196216 106224 196222 106276
rect 197630 106264 197636 106276
rect 197591 106236 197636 106264
rect 197630 106224 197636 106236
rect 197688 106224 197694 106276
rect 200298 106224 200304 106276
rect 200356 106224 200362 106276
rect 218238 106224 218244 106276
rect 218296 106224 218302 106276
rect 220998 106224 221004 106276
rect 221056 106224 221062 106276
rect 222473 106267 222531 106273
rect 222473 106233 222485 106267
rect 222519 106264 222531 106267
rect 222562 106264 222568 106276
rect 222519 106236 222568 106264
rect 222519 106233 222531 106236
rect 222473 106227 222531 106233
rect 222562 106224 222568 106236
rect 222620 106224 222626 106276
rect 238754 106224 238760 106276
rect 238812 106264 238818 106276
rect 239030 106264 239036 106276
rect 238812 106236 239036 106264
rect 238812 106224 238818 106236
rect 239030 106224 239036 106236
rect 239088 106224 239094 106276
rect 240410 106264 240416 106276
rect 240371 106236 240416 106264
rect 240410 106224 240416 106236
rect 240468 106224 240474 106276
rect 200316 106140 200344 106224
rect 200298 106088 200304 106140
rect 200356 106088 200362 106140
rect 219618 104932 219624 104984
rect 219676 104932 219682 104984
rect 180981 104907 181039 104913
rect 180981 104873 180993 104907
rect 181027 104904 181039 104907
rect 181162 104904 181168 104916
rect 181027 104876 181168 104904
rect 181027 104873 181039 104876
rect 180981 104867 181039 104873
rect 181162 104864 181168 104876
rect 181220 104864 181226 104916
rect 182450 104904 182456 104916
rect 182411 104876 182456 104904
rect 182450 104864 182456 104876
rect 182508 104864 182514 104916
rect 183830 104864 183836 104916
rect 183888 104904 183894 104916
rect 183922 104904 183928 104916
rect 183888 104876 183928 104904
rect 183888 104864 183894 104876
rect 183922 104864 183928 104876
rect 183980 104864 183986 104916
rect 174170 104836 174176 104848
rect 174131 104808 174176 104836
rect 174170 104796 174176 104808
rect 174228 104796 174234 104848
rect 219636 104780 219664 104932
rect 385034 104796 385040 104848
rect 385092 104836 385098 104848
rect 385092 104808 385137 104836
rect 385092 104796 385098 104808
rect 218238 104768 218244 104780
rect 218199 104740 218244 104768
rect 218238 104728 218244 104740
rect 218296 104728 218302 104780
rect 219618 104728 219624 104780
rect 219676 104728 219682 104780
rect 182358 103572 182364 103624
rect 182416 103612 182422 103624
rect 182453 103615 182511 103621
rect 182453 103612 182465 103615
rect 182416 103584 182465 103612
rect 182416 103572 182422 103584
rect 182453 103581 182465 103584
rect 182499 103581 182511 103615
rect 182453 103575 182511 103581
rect 158901 103547 158959 103553
rect 158901 103513 158913 103547
rect 158947 103544 158959 103547
rect 159082 103544 159088 103556
rect 158947 103516 159088 103544
rect 158947 103513 158959 103516
rect 158901 103507 158959 103513
rect 159082 103504 159088 103516
rect 159140 103504 159146 103556
rect 223850 103544 223856 103556
rect 223776 103516 223856 103544
rect 223776 103408 223804 103516
rect 223850 103504 223856 103516
rect 223908 103504 223914 103556
rect 223942 103408 223948 103420
rect 223776 103380 223948 103408
rect 223942 103368 223948 103380
rect 224000 103368 224006 103420
rect 182450 102076 182456 102128
rect 182508 102116 182514 102128
rect 182545 102119 182603 102125
rect 182545 102116 182557 102119
rect 182508 102088 182557 102116
rect 182508 102076 182514 102088
rect 182545 102085 182557 102088
rect 182591 102085 182603 102119
rect 182545 102079 182603 102085
rect 183830 101396 183836 101448
rect 183888 101396 183894 101448
rect 239030 101396 239036 101448
rect 239088 101396 239094 101448
rect 183848 101312 183876 101396
rect 239048 101312 239076 101396
rect 183830 101260 183836 101312
rect 183888 101260 183894 101312
rect 239030 101260 239036 101312
rect 239088 101260 239094 101312
rect 218238 100008 218244 100020
rect 218199 99980 218244 100008
rect 218238 99968 218244 99980
rect 218296 99968 218302 100020
rect 217042 99464 217048 99476
rect 217003 99436 217048 99464
rect 217042 99424 217048 99436
rect 217100 99424 217106 99476
rect 157518 99356 157524 99408
rect 157576 99396 157582 99408
rect 157702 99396 157708 99408
rect 157576 99368 157708 99396
rect 157576 99356 157582 99368
rect 157702 99356 157708 99368
rect 157760 99356 157766 99408
rect 163038 99356 163044 99408
rect 163096 99396 163102 99408
rect 163222 99396 163228 99408
rect 163096 99368 163228 99396
rect 163096 99356 163102 99368
rect 163222 99356 163228 99368
rect 163280 99356 163286 99408
rect 181070 99356 181076 99408
rect 181128 99396 181134 99408
rect 181128 99368 181208 99396
rect 181128 99356 181134 99368
rect 181180 99340 181208 99368
rect 205818 99356 205824 99408
rect 205876 99356 205882 99408
rect 207290 99356 207296 99408
rect 207348 99356 207354 99408
rect 181162 99288 181168 99340
rect 181220 99288 181226 99340
rect 205836 99328 205864 99356
rect 205910 99328 205916 99340
rect 205836 99300 205916 99328
rect 205910 99288 205916 99300
rect 205968 99288 205974 99340
rect 207308 99328 207336 99356
rect 207382 99328 207388 99340
rect 207308 99300 207388 99328
rect 207382 99288 207388 99300
rect 207440 99288 207446 99340
rect 219529 98719 219587 98725
rect 219529 98685 219541 98719
rect 219575 98716 219587 98719
rect 219618 98716 219624 98728
rect 219575 98688 219624 98716
rect 219575 98685 219587 98688
rect 219529 98679 219587 98685
rect 219618 98676 219624 98688
rect 219676 98676 219682 98728
rect 256694 97928 256700 97980
rect 256752 97968 256758 97980
rect 256878 97968 256884 97980
rect 256752 97940 256884 97968
rect 256752 97928 256758 97940
rect 256878 97928 256884 97940
rect 256936 97928 256942 97980
rect 182450 97248 182456 97300
rect 182508 97288 182514 97300
rect 182545 97291 182603 97297
rect 182545 97288 182557 97291
rect 182508 97260 182557 97288
rect 182508 97248 182514 97260
rect 182545 97257 182557 97260
rect 182591 97257 182603 97291
rect 182545 97251 182603 97257
rect 196158 96676 196164 96688
rect 196119 96648 196164 96676
rect 196158 96636 196164 96648
rect 196216 96636 196222 96688
rect 197630 96676 197636 96688
rect 197591 96648 197636 96676
rect 197630 96636 197636 96648
rect 197688 96636 197694 96688
rect 222470 96676 222476 96688
rect 222431 96648 222476 96676
rect 222470 96636 222476 96648
rect 222528 96636 222534 96688
rect 240410 96676 240416 96688
rect 240371 96648 240416 96676
rect 240410 96636 240416 96648
rect 240468 96636 240474 96688
rect 163130 96608 163136 96620
rect 163091 96580 163136 96608
rect 163130 96568 163136 96580
rect 163188 96568 163194 96620
rect 185026 96568 185032 96620
rect 185084 96608 185090 96620
rect 185210 96608 185216 96620
rect 185084 96580 185216 96608
rect 185084 96568 185090 96580
rect 185210 96568 185216 96580
rect 185268 96568 185274 96620
rect 217042 96608 217048 96620
rect 217003 96580 217048 96608
rect 217042 96568 217048 96580
rect 217100 96568 217106 96620
rect 158898 95208 158904 95260
rect 158956 95248 158962 95260
rect 159082 95248 159088 95260
rect 158956 95220 159088 95248
rect 158956 95208 158962 95220
rect 159082 95208 159088 95220
rect 159140 95208 159146 95260
rect 168558 95208 168564 95260
rect 168616 95248 168622 95260
rect 168650 95248 168656 95260
rect 168616 95220 168656 95248
rect 168616 95208 168622 95220
rect 168650 95208 168656 95220
rect 168708 95208 168714 95260
rect 174173 95251 174231 95257
rect 174173 95217 174185 95251
rect 174219 95248 174231 95251
rect 174262 95248 174268 95260
rect 174219 95220 174268 95248
rect 174219 95217 174231 95220
rect 174173 95211 174231 95217
rect 174262 95208 174268 95220
rect 174320 95208 174326 95260
rect 181070 95180 181076 95192
rect 181031 95152 181076 95180
rect 181070 95140 181076 95152
rect 181128 95140 181134 95192
rect 185026 95180 185032 95192
rect 184987 95152 185032 95180
rect 185026 95140 185032 95152
rect 185084 95140 185090 95192
rect 218238 95180 218244 95192
rect 218199 95152 218244 95180
rect 218238 95140 218244 95152
rect 218296 95140 218302 95192
rect 158898 95112 158904 95124
rect 158859 95084 158904 95112
rect 158898 95072 158904 95084
rect 158956 95072 158962 95124
rect 378134 93848 378140 93900
rect 378192 93888 378198 93900
rect 378318 93888 378324 93900
rect 378192 93860 378324 93888
rect 378192 93848 378198 93860
rect 378318 93848 378324 93860
rect 378376 93848 378382 93900
rect 385037 93891 385095 93897
rect 385037 93857 385049 93891
rect 385083 93888 385095 93891
rect 385126 93888 385132 93900
rect 385083 93860 385132 93888
rect 385083 93857 385095 93860
rect 385037 93851 385095 93857
rect 385126 93848 385132 93860
rect 385184 93848 385190 93900
rect 3602 93780 3608 93832
rect 3660 93820 3666 93832
rect 152734 93820 152740 93832
rect 3660 93792 152740 93820
rect 3660 93780 3666 93792
rect 152734 93780 152740 93792
rect 152792 93780 152798 93832
rect 219437 92463 219495 92469
rect 219437 92429 219449 92463
rect 219483 92460 219495 92463
rect 219529 92463 219587 92469
rect 219529 92460 219541 92463
rect 219483 92432 219541 92460
rect 219483 92429 219495 92432
rect 219437 92423 219495 92429
rect 219529 92429 219541 92432
rect 219575 92429 219587 92463
rect 227990 92460 227996 92472
rect 227951 92432 227996 92460
rect 219529 92423 219587 92429
rect 227990 92420 227996 92432
rect 228048 92420 228054 92472
rect 218241 91851 218299 91857
rect 218241 91817 218253 91851
rect 218287 91848 218299 91851
rect 218330 91848 218336 91860
rect 218287 91820 218336 91848
rect 218287 91817 218299 91820
rect 218241 91811 218299 91817
rect 218330 91808 218336 91820
rect 218388 91808 218394 91860
rect 156230 89700 156236 89752
rect 156288 89740 156294 89752
rect 156414 89740 156420 89752
rect 156288 89712 156420 89740
rect 156288 89700 156294 89712
rect 156414 89700 156420 89712
rect 156472 89700 156478 89752
rect 157610 89700 157616 89752
rect 157668 89700 157674 89752
rect 174078 89700 174084 89752
rect 174136 89740 174142 89752
rect 174262 89740 174268 89752
rect 174136 89712 174268 89740
rect 174136 89700 174142 89712
rect 174262 89700 174268 89712
rect 174320 89700 174326 89752
rect 193398 89700 193404 89752
rect 193456 89740 193462 89752
rect 193582 89740 193588 89752
rect 193456 89712 193588 89740
rect 193456 89700 193462 89712
rect 193582 89700 193588 89712
rect 193640 89700 193646 89752
rect 205726 89700 205732 89752
rect 205784 89740 205790 89752
rect 205910 89740 205916 89752
rect 205784 89712 205916 89740
rect 205784 89700 205790 89712
rect 205910 89700 205916 89712
rect 205968 89700 205974 89752
rect 157628 89604 157656 89700
rect 163130 89672 163136 89684
rect 163091 89644 163136 89672
rect 163130 89632 163136 89644
rect 163188 89632 163194 89684
rect 157702 89604 157708 89616
rect 157628 89576 157708 89604
rect 157702 89564 157708 89576
rect 157760 89564 157766 89616
rect 392854 88272 392860 88324
rect 392912 88312 392918 88324
rect 579890 88312 579896 88324
rect 392912 88284 579896 88312
rect 392912 88272 392918 88284
rect 579890 88272 579896 88284
rect 579948 88272 579954 88324
rect 200298 86912 200304 86964
rect 200356 86912 200362 86964
rect 209869 86955 209927 86961
rect 209869 86921 209881 86955
rect 209915 86952 209927 86955
rect 209958 86952 209964 86964
rect 209915 86924 209964 86952
rect 209915 86921 209927 86924
rect 209869 86915 209927 86921
rect 209958 86912 209964 86924
rect 210016 86912 210022 86964
rect 216950 86912 216956 86964
rect 217008 86952 217014 86964
rect 217042 86952 217048 86964
rect 217008 86924 217048 86952
rect 217008 86912 217014 86924
rect 217042 86912 217048 86924
rect 217100 86912 217106 86964
rect 239030 86952 239036 86964
rect 238991 86924 239036 86952
rect 239030 86912 239036 86924
rect 239088 86912 239094 86964
rect 240410 86952 240416 86964
rect 240371 86924 240416 86952
rect 240410 86912 240416 86924
rect 240468 86912 240474 86964
rect 200316 86828 200344 86912
rect 200298 86776 200304 86828
rect 200356 86776 200362 86828
rect 183830 85796 183836 85808
rect 183791 85768 183836 85796
rect 183830 85756 183836 85768
rect 183888 85756 183894 85808
rect 158901 85595 158959 85601
rect 158901 85561 158913 85595
rect 158947 85592 158959 85595
rect 158990 85592 158996 85604
rect 158947 85564 158996 85592
rect 158947 85561 158959 85564
rect 158901 85555 158959 85561
rect 158990 85552 158996 85564
rect 159048 85552 159054 85604
rect 181073 85595 181131 85601
rect 181073 85561 181085 85595
rect 181119 85592 181131 85595
rect 181162 85592 181168 85604
rect 181119 85564 181168 85592
rect 181119 85561 181131 85564
rect 181073 85555 181131 85561
rect 181162 85552 181168 85564
rect 181220 85552 181226 85604
rect 185029 85595 185087 85601
rect 185029 85561 185041 85595
rect 185075 85592 185087 85595
rect 185210 85592 185216 85604
rect 185075 85564 185216 85592
rect 185075 85561 185087 85564
rect 185029 85555 185087 85561
rect 185210 85552 185216 85564
rect 185268 85552 185274 85604
rect 220998 85552 221004 85604
rect 221056 85592 221062 85604
rect 221090 85592 221096 85604
rect 221056 85564 221096 85592
rect 221056 85552 221062 85564
rect 221090 85552 221096 85564
rect 221148 85552 221154 85604
rect 223850 85552 223856 85604
rect 223908 85592 223914 85604
rect 223942 85592 223948 85604
rect 223908 85564 223948 85592
rect 223908 85552 223914 85564
rect 223942 85552 223948 85564
rect 224000 85552 224006 85604
rect 174170 85524 174176 85536
rect 174131 85496 174176 85524
rect 174170 85484 174176 85496
rect 174228 85484 174234 85536
rect 183830 84232 183836 84244
rect 183791 84204 183836 84232
rect 183830 84192 183836 84204
rect 183888 84192 183894 84244
rect 182450 84164 182456 84176
rect 182411 84136 182456 84164
rect 182450 84124 182456 84136
rect 182508 84124 182514 84176
rect 385037 84167 385095 84173
rect 385037 84133 385049 84167
rect 385083 84164 385095 84167
rect 385126 84164 385132 84176
rect 385083 84136 385132 84164
rect 385083 84133 385095 84136
rect 385037 84127 385095 84133
rect 385126 84124 385132 84136
rect 385184 84124 385190 84176
rect 219437 82875 219495 82881
rect 219437 82841 219449 82875
rect 219483 82872 219495 82875
rect 219621 82875 219679 82881
rect 219621 82872 219633 82875
rect 219483 82844 219633 82872
rect 219483 82841 219495 82844
rect 219437 82835 219495 82841
rect 219621 82841 219633 82844
rect 219667 82841 219679 82875
rect 219621 82835 219679 82841
rect 227993 82875 228051 82881
rect 227993 82841 228005 82875
rect 228039 82872 228051 82875
rect 228082 82872 228088 82884
rect 228039 82844 228088 82872
rect 228039 82841 228051 82844
rect 227993 82835 228051 82841
rect 228082 82832 228088 82844
rect 228140 82832 228146 82884
rect 207198 80152 207204 80164
rect 207124 80124 207204 80152
rect 157518 80044 157524 80096
rect 157576 80084 157582 80096
rect 157702 80084 157708 80096
rect 157576 80056 157708 80084
rect 157576 80044 157582 80056
rect 157702 80044 157708 80056
rect 157760 80044 157766 80096
rect 163038 80044 163044 80096
rect 163096 80084 163102 80096
rect 163222 80084 163228 80096
rect 163096 80056 163228 80084
rect 163096 80044 163102 80056
rect 163222 80044 163228 80056
rect 163280 80044 163286 80096
rect 181070 80044 181076 80096
rect 181128 80044 181134 80096
rect 205818 80044 205824 80096
rect 205876 80044 205882 80096
rect 3050 79976 3056 80028
rect 3108 80016 3114 80028
rect 152826 80016 152832 80028
rect 3108 79988 152832 80016
rect 3108 79976 3114 79988
rect 152826 79976 152832 79988
rect 152884 79976 152890 80028
rect 181088 80016 181116 80044
rect 181162 80016 181168 80028
rect 181088 79988 181168 80016
rect 181162 79976 181168 79988
rect 181220 79976 181226 80028
rect 205836 79948 205864 80044
rect 207124 80028 207152 80124
rect 207198 80112 207204 80124
rect 207256 80112 207262 80164
rect 256878 80044 256884 80096
rect 256936 80044 256942 80096
rect 207106 79976 207112 80028
rect 207164 79976 207170 80028
rect 205910 79948 205916 79960
rect 205836 79920 205916 79948
rect 205910 79908 205916 79920
rect 205968 79908 205974 79960
rect 256896 79948 256924 80044
rect 256970 79948 256976 79960
rect 256896 79920 256976 79948
rect 256970 79908 256976 79920
rect 257028 79908 257034 79960
rect 182450 79336 182456 79348
rect 182411 79308 182456 79336
rect 182450 79296 182456 79308
rect 182508 79296 182514 79348
rect 227993 77979 228051 77985
rect 227993 77945 228005 77979
rect 228039 77976 228051 77979
rect 228082 77976 228088 77988
rect 228039 77948 228088 77976
rect 228039 77945 228051 77948
rect 227993 77939 228051 77945
rect 228082 77936 228088 77948
rect 228140 77936 228146 77988
rect 222562 77364 222568 77376
rect 222488 77336 222568 77364
rect 222488 77308 222516 77336
rect 222562 77324 222568 77336
rect 222620 77324 222626 77376
rect 209866 77296 209872 77308
rect 209827 77268 209872 77296
rect 209866 77256 209872 77268
rect 209924 77256 209930 77308
rect 222470 77256 222476 77308
rect 222528 77256 222534 77308
rect 239030 77296 239036 77308
rect 238991 77268 239036 77296
rect 239030 77256 239036 77268
rect 239088 77256 239094 77308
rect 240410 77296 240416 77308
rect 240371 77268 240416 77296
rect 240410 77256 240416 77268
rect 240468 77256 240474 77308
rect 207106 77228 207112 77240
rect 207067 77200 207112 77228
rect 207106 77188 207112 77200
rect 207164 77188 207170 77240
rect 256881 77231 256939 77237
rect 256881 77197 256893 77231
rect 256927 77228 256939 77231
rect 256970 77228 256976 77240
rect 256927 77200 256976 77228
rect 256927 77197 256939 77200
rect 256881 77191 256939 77197
rect 256970 77188 256976 77200
rect 257028 77188 257034 77240
rect 392762 77188 392768 77240
rect 392820 77228 392826 77240
rect 579890 77228 579896 77240
rect 392820 77200 579896 77228
rect 392820 77188 392826 77200
rect 579890 77188 579896 77200
rect 579948 77188 579954 77240
rect 158714 75896 158720 75948
rect 158772 75936 158778 75948
rect 158898 75936 158904 75948
rect 158772 75908 158904 75936
rect 158772 75896 158778 75908
rect 158898 75896 158904 75908
rect 158956 75896 158962 75948
rect 174173 75939 174231 75945
rect 174173 75905 174185 75939
rect 174219 75936 174231 75939
rect 174262 75936 174268 75948
rect 174219 75908 174268 75936
rect 174219 75905 174231 75908
rect 174173 75899 174231 75905
rect 174262 75896 174268 75908
rect 174320 75896 174326 75948
rect 218238 75896 218244 75948
rect 218296 75936 218302 75948
rect 218330 75936 218336 75948
rect 218296 75908 218336 75936
rect 218296 75896 218302 75908
rect 218330 75896 218336 75908
rect 218388 75896 218394 75948
rect 219618 75936 219624 75948
rect 219579 75908 219624 75936
rect 219618 75896 219624 75908
rect 219676 75896 219682 75948
rect 181070 75868 181076 75880
rect 181031 75840 181076 75868
rect 181070 75828 181076 75840
rect 181128 75828 181134 75880
rect 378134 74536 378140 74588
rect 378192 74576 378198 74588
rect 378318 74576 378324 74588
rect 378192 74548 378324 74576
rect 378192 74536 378198 74548
rect 378318 74536 378324 74548
rect 378376 74536 378382 74588
rect 222470 73148 222476 73160
rect 222431 73120 222476 73148
rect 222470 73108 222476 73120
rect 222528 73108 222534 73160
rect 183830 70700 183836 70712
rect 183791 70672 183836 70700
rect 183830 70660 183836 70672
rect 183888 70660 183894 70712
rect 157610 70388 157616 70440
rect 157668 70388 157674 70440
rect 163130 70388 163136 70440
rect 163188 70388 163194 70440
rect 185118 70388 185124 70440
rect 185176 70388 185182 70440
rect 157628 70292 157656 70388
rect 157702 70292 157708 70304
rect 157628 70264 157708 70292
rect 157702 70252 157708 70264
rect 157760 70252 157766 70304
rect 163148 70292 163176 70388
rect 163222 70292 163228 70304
rect 163148 70264 163228 70292
rect 163222 70252 163228 70264
rect 163280 70252 163286 70304
rect 185136 70292 185164 70388
rect 207109 70363 207167 70369
rect 207109 70329 207121 70363
rect 207155 70360 207167 70363
rect 207198 70360 207204 70372
rect 207155 70332 207204 70360
rect 207155 70329 207167 70332
rect 207109 70323 207167 70329
rect 207198 70320 207204 70332
rect 207256 70320 207262 70372
rect 185210 70292 185216 70304
rect 185136 70264 185216 70292
rect 185210 70252 185216 70264
rect 185268 70252 185274 70304
rect 205910 67708 205916 67720
rect 205836 67680 205916 67708
rect 205836 67652 205864 67680
rect 205910 67668 205916 67680
rect 205968 67668 205974 67720
rect 168558 67600 168564 67652
rect 168616 67640 168622 67652
rect 168650 67640 168656 67652
rect 168616 67612 168656 67640
rect 168616 67600 168622 67612
rect 168650 67600 168656 67612
rect 168708 67600 168714 67652
rect 205818 67600 205824 67652
rect 205876 67600 205882 67652
rect 256878 67640 256884 67652
rect 256839 67612 256884 67640
rect 256878 67600 256884 67612
rect 256936 67600 256942 67652
rect 216953 67575 217011 67581
rect 216953 67541 216965 67575
rect 216999 67572 217011 67575
rect 217042 67572 217048 67584
rect 216999 67544 217048 67572
rect 216999 67541 217011 67544
rect 216953 67535 217011 67541
rect 217042 67532 217048 67544
rect 217100 67532 217106 67584
rect 240410 67572 240416 67584
rect 240371 67544 240416 67572
rect 240410 67532 240416 67544
rect 240468 67532 240474 67584
rect 221090 66348 221096 66360
rect 221016 66320 221096 66348
rect 221016 66292 221044 66320
rect 221090 66308 221096 66320
rect 221148 66308 221154 66360
rect 225322 66348 225328 66360
rect 225248 66320 225328 66348
rect 225248 66292 225276 66320
rect 225322 66308 225328 66320
rect 225380 66308 225386 66360
rect 226702 66348 226708 66360
rect 226628 66320 226708 66348
rect 226628 66292 226656 66320
rect 226702 66308 226708 66320
rect 226760 66308 226766 66360
rect 174170 66240 174176 66292
rect 174228 66280 174234 66292
rect 174262 66280 174268 66292
rect 174228 66252 174268 66280
rect 174228 66240 174234 66252
rect 174262 66240 174268 66252
rect 174320 66240 174326 66292
rect 181073 66283 181131 66289
rect 181073 66249 181085 66283
rect 181119 66280 181131 66283
rect 181162 66280 181168 66292
rect 181119 66252 181168 66280
rect 181119 66249 181131 66252
rect 181073 66243 181131 66249
rect 181162 66240 181168 66252
rect 181220 66240 181226 66292
rect 182358 66240 182364 66292
rect 182416 66280 182422 66292
rect 182450 66280 182456 66292
rect 182416 66252 182456 66280
rect 182416 66240 182422 66252
rect 182450 66240 182456 66252
rect 182508 66240 182514 66292
rect 183830 66280 183836 66292
rect 183791 66252 183836 66280
rect 183830 66240 183836 66252
rect 183888 66240 183894 66292
rect 220998 66240 221004 66292
rect 221056 66240 221062 66292
rect 225230 66240 225236 66292
rect 225288 66240 225294 66292
rect 226610 66240 226616 66292
rect 226668 66240 226674 66292
rect 385034 66240 385040 66292
rect 385092 66280 385098 66292
rect 385092 66252 385137 66280
rect 385092 66240 385098 66252
rect 158990 66212 158996 66224
rect 158951 66184 158996 66212
rect 158990 66172 158996 66184
rect 159048 66172 159054 66224
rect 237282 66212 237288 66224
rect 237243 66184 237288 66212
rect 237282 66172 237288 66184
rect 237340 66172 237346 66224
rect 238662 66212 238668 66224
rect 238623 66184 238668 66212
rect 238662 66172 238668 66184
rect 238720 66172 238726 66224
rect 223758 64880 223764 64932
rect 223816 64920 223822 64932
rect 223850 64920 223856 64932
rect 223816 64892 223856 64920
rect 223816 64880 223822 64892
rect 223850 64880 223856 64892
rect 223908 64880 223914 64932
rect 227990 64920 227996 64932
rect 227951 64892 227996 64920
rect 227990 64880 227996 64892
rect 228048 64880 228054 64932
rect 182358 64852 182364 64864
rect 182319 64824 182364 64852
rect 182358 64812 182364 64824
rect 182416 64812 182422 64864
rect 183830 64852 183836 64864
rect 183791 64824 183836 64852
rect 183830 64812 183836 64824
rect 183888 64812 183894 64864
rect 185210 64852 185216 64864
rect 185171 64824 185216 64852
rect 185210 64812 185216 64824
rect 185268 64812 185274 64864
rect 393958 64812 393964 64864
rect 394016 64852 394022 64864
rect 580166 64852 580172 64864
rect 394016 64824 580172 64852
rect 394016 64812 394022 64824
rect 580166 64812 580172 64824
rect 580224 64812 580230 64864
rect 222473 63563 222531 63569
rect 222473 63529 222485 63563
rect 222519 63560 222531 63563
rect 222654 63560 222660 63572
rect 222519 63532 222660 63560
rect 222519 63529 222531 63532
rect 222473 63523 222531 63529
rect 222654 63520 222660 63532
rect 222712 63520 222718 63572
rect 240410 62744 240416 62756
rect 240371 62716 240416 62744
rect 240410 62704 240416 62716
rect 240468 62704 240474 62756
rect 180981 60843 181039 60849
rect 180981 60809 180993 60843
rect 181027 60840 181039 60843
rect 181162 60840 181168 60852
rect 181027 60812 181168 60840
rect 181027 60809 181039 60812
rect 180981 60803 181039 60809
rect 181162 60800 181168 60812
rect 181220 60800 181226 60852
rect 207198 60664 207204 60716
rect 207256 60704 207262 60716
rect 207382 60704 207388 60716
rect 207256 60676 207388 60704
rect 207256 60664 207262 60676
rect 207382 60664 207388 60676
rect 207440 60664 207446 60716
rect 209958 60664 209964 60716
rect 210016 60704 210022 60716
rect 210142 60704 210148 60716
rect 210016 60676 210148 60704
rect 210016 60664 210022 60676
rect 210142 60664 210148 60676
rect 210200 60664 210206 60716
rect 185118 59168 185124 59220
rect 185176 59208 185182 59220
rect 185213 59211 185271 59217
rect 185213 59208 185225 59211
rect 185176 59180 185225 59208
rect 185176 59168 185182 59180
rect 185213 59177 185225 59180
rect 185259 59177 185271 59211
rect 185213 59171 185271 59177
rect 223758 58012 223764 58064
rect 223816 58012 223822 58064
rect 168558 57944 168564 57996
rect 168616 57984 168622 57996
rect 168650 57984 168656 57996
rect 168616 57956 168656 57984
rect 168616 57944 168622 57956
rect 168650 57944 168656 57956
rect 168708 57944 168714 57996
rect 219526 57944 219532 57996
rect 219584 57984 219590 57996
rect 219618 57984 219624 57996
rect 219584 57956 219624 57984
rect 219584 57944 219590 57956
rect 219618 57944 219624 57956
rect 219676 57944 219682 57996
rect 220998 57944 221004 57996
rect 221056 57984 221062 57996
rect 221090 57984 221096 57996
rect 221056 57956 221096 57984
rect 221056 57944 221062 57956
rect 221090 57944 221096 57956
rect 221148 57944 221154 57996
rect 223776 57928 223804 58012
rect 225230 57944 225236 57996
rect 225288 57984 225294 57996
rect 225322 57984 225328 57996
rect 225288 57956 225328 57984
rect 225288 57944 225294 57956
rect 225322 57944 225328 57956
rect 225380 57944 225386 57996
rect 256694 57944 256700 57996
rect 256752 57984 256758 57996
rect 256970 57984 256976 57996
rect 256752 57956 256976 57984
rect 256752 57944 256758 57956
rect 256970 57944 256976 57956
rect 257028 57944 257034 57996
rect 180978 57916 180984 57928
rect 180939 57888 180984 57916
rect 180978 57876 180984 57888
rect 181036 57876 181042 57928
rect 193493 57919 193551 57925
rect 193493 57885 193505 57919
rect 193539 57916 193551 57919
rect 193582 57916 193588 57928
rect 193539 57888 193588 57916
rect 193539 57885 193551 57888
rect 193493 57879 193551 57885
rect 193582 57876 193588 57888
rect 193640 57876 193646 57928
rect 210053 57919 210111 57925
rect 210053 57885 210065 57919
rect 210099 57916 210111 57919
rect 210142 57916 210148 57928
rect 210099 57888 210148 57916
rect 210099 57885 210111 57888
rect 210053 57879 210111 57885
rect 210142 57876 210148 57888
rect 210200 57876 210206 57928
rect 223758 57876 223764 57928
rect 223816 57876 223822 57928
rect 239030 57916 239036 57928
rect 238991 57888 239036 57916
rect 239030 57876 239036 57888
rect 239088 57876 239094 57928
rect 158990 56624 158996 56636
rect 158951 56596 158996 56624
rect 158990 56584 158996 56596
rect 159048 56584 159054 56636
rect 216953 56627 217011 56633
rect 216953 56593 216965 56627
rect 216999 56624 217011 56627
rect 217042 56624 217048 56636
rect 216999 56596 217048 56624
rect 216999 56593 217011 56596
rect 216953 56587 217011 56593
rect 217042 56584 217048 56596
rect 217100 56584 217106 56636
rect 237282 56624 237288 56636
rect 237243 56596 237288 56624
rect 237282 56584 237288 56596
rect 237340 56584 237346 56636
rect 238662 56624 238668 56636
rect 238623 56596 238668 56624
rect 238662 56584 238668 56596
rect 238720 56584 238726 56636
rect 180978 56556 180984 56568
rect 180939 56528 180984 56556
rect 180978 56516 180984 56528
rect 181036 56516 181042 56568
rect 218241 56559 218299 56565
rect 218241 56525 218253 56559
rect 218287 56556 218299 56559
rect 218330 56556 218336 56568
rect 218287 56528 218336 56556
rect 218287 56525 218299 56528
rect 218241 56519 218299 56525
rect 218330 56516 218336 56528
rect 218388 56516 218394 56568
rect 183830 55264 183836 55276
rect 183791 55236 183836 55264
rect 183830 55224 183836 55236
rect 183888 55224 183894 55276
rect 378134 55224 378140 55276
rect 378192 55264 378198 55276
rect 378318 55264 378324 55276
rect 378192 55236 378324 55264
rect 378192 55224 378198 55236
rect 378318 55224 378324 55236
rect 378376 55224 378382 55276
rect 222565 54655 222623 54661
rect 222565 54621 222577 54655
rect 222611 54652 222623 54655
rect 222654 54652 222660 54664
rect 222611 54624 222660 54652
rect 222611 54621 222623 54624
rect 222565 54615 222623 54621
rect 222654 54612 222660 54624
rect 222712 54612 222718 54664
rect 207382 51116 207388 51128
rect 207308 51088 207388 51116
rect 207308 51060 207336 51088
rect 207382 51076 207388 51088
rect 207440 51076 207446 51128
rect 3050 51008 3056 51060
rect 3108 51048 3114 51060
rect 152550 51048 152556 51060
rect 3108 51020 152556 51048
rect 3108 51008 3114 51020
rect 152550 51008 152556 51020
rect 152608 51008 152614 51060
rect 207290 51008 207296 51060
rect 207348 51008 207354 51060
rect 385126 51008 385132 51060
rect 385184 51048 385190 51060
rect 385310 51048 385316 51060
rect 385184 51020 385316 51048
rect 385184 51008 385190 51020
rect 385310 51008 385316 51020
rect 385368 51008 385374 51060
rect 205910 48396 205916 48408
rect 205836 48368 205916 48396
rect 205836 48340 205864 48368
rect 205910 48356 205916 48368
rect 205968 48356 205974 48408
rect 219618 48396 219624 48408
rect 219544 48368 219624 48396
rect 219544 48340 219572 48368
rect 219618 48356 219624 48368
rect 219676 48356 219682 48408
rect 221090 48396 221096 48408
rect 221016 48368 221096 48396
rect 221016 48340 221044 48368
rect 221090 48356 221096 48368
rect 221148 48356 221154 48408
rect 158990 48328 158996 48340
rect 158916 48300 158996 48328
rect 158916 48272 158944 48300
rect 158990 48288 158996 48300
rect 159048 48288 159054 48340
rect 182358 48328 182364 48340
rect 182319 48300 182364 48328
rect 182358 48288 182364 48300
rect 182416 48288 182422 48340
rect 193490 48328 193496 48340
rect 193451 48300 193496 48328
rect 193490 48288 193496 48300
rect 193548 48288 193554 48340
rect 205818 48288 205824 48340
rect 205876 48288 205882 48340
rect 210050 48328 210056 48340
rect 210011 48300 210056 48328
rect 210050 48288 210056 48300
rect 210108 48288 210114 48340
rect 219526 48288 219532 48340
rect 219584 48288 219590 48340
rect 220998 48288 221004 48340
rect 221056 48288 221062 48340
rect 237190 48288 237196 48340
rect 237248 48328 237254 48340
rect 237282 48328 237288 48340
rect 237248 48300 237288 48328
rect 237248 48288 237254 48300
rect 237282 48288 237288 48300
rect 237340 48288 237346 48340
rect 238662 48288 238668 48340
rect 238720 48328 238726 48340
rect 238754 48328 238760 48340
rect 238720 48300 238760 48328
rect 238720 48288 238726 48300
rect 238754 48288 238760 48300
rect 238812 48288 238818 48340
rect 239030 48328 239036 48340
rect 238991 48300 239036 48328
rect 239030 48288 239036 48300
rect 239088 48288 239094 48340
rect 256510 48288 256516 48340
rect 256568 48328 256574 48340
rect 256878 48328 256884 48340
rect 256568 48300 256884 48328
rect 256568 48288 256574 48300
rect 256878 48288 256884 48300
rect 256936 48288 256942 48340
rect 158898 48220 158904 48272
rect 158956 48220 158962 48272
rect 223758 48220 223764 48272
rect 223816 48260 223822 48272
rect 223942 48260 223948 48272
rect 223816 48232 223948 48260
rect 223816 48220 223822 48232
rect 223942 48220 223948 48232
rect 224000 48220 224006 48272
rect 225230 48220 225236 48272
rect 225288 48260 225294 48272
rect 225414 48260 225420 48272
rect 225288 48232 225420 48260
rect 225288 48220 225294 48232
rect 225414 48220 225420 48232
rect 225472 48220 225478 48272
rect 180981 46971 181039 46977
rect 180981 46937 180993 46971
rect 181027 46968 181039 46971
rect 181162 46968 181168 46980
rect 181027 46940 181168 46968
rect 181027 46937 181039 46940
rect 180981 46931 181039 46937
rect 181162 46928 181168 46940
rect 181220 46928 181226 46980
rect 218238 46968 218244 46980
rect 218199 46940 218244 46968
rect 218238 46928 218244 46940
rect 218296 46928 218302 46980
rect 158898 46900 158904 46912
rect 158859 46872 158904 46900
rect 158898 46860 158904 46872
rect 158956 46860 158962 46912
rect 182358 46900 182364 46912
rect 182319 46872 182364 46900
rect 182358 46860 182364 46872
rect 182416 46860 182422 46912
rect 210050 46900 210056 46912
rect 210011 46872 210056 46900
rect 210050 46860 210056 46872
rect 210108 46860 210114 46912
rect 220998 46900 221004 46912
rect 220959 46872 221004 46900
rect 220998 46860 221004 46872
rect 221056 46860 221062 46912
rect 226610 46860 226616 46912
rect 226668 46900 226674 46912
rect 226702 46900 226708 46912
rect 226668 46872 226708 46900
rect 226668 46860 226674 46872
rect 226702 46860 226708 46872
rect 226760 46860 226766 46912
rect 237282 46900 237288 46912
rect 237243 46872 237288 46900
rect 237282 46860 237288 46872
rect 237340 46860 237346 46912
rect 238662 46900 238668 46912
rect 238623 46872 238668 46900
rect 238662 46860 238668 46872
rect 238720 46860 238726 46912
rect 183922 45568 183928 45620
rect 183980 45608 183986 45620
rect 184014 45608 184020 45620
rect 183980 45580 184020 45608
rect 183980 45568 183986 45580
rect 184014 45568 184020 45580
rect 184072 45568 184078 45620
rect 222562 45608 222568 45620
rect 222523 45580 222568 45608
rect 222562 45568 222568 45580
rect 222620 45568 222626 45620
rect 185118 45500 185124 45552
rect 185176 45540 185182 45552
rect 185394 45540 185400 45552
rect 185176 45512 185400 45540
rect 185176 45500 185182 45512
rect 185394 45500 185400 45512
rect 185452 45500 185458 45552
rect 181162 41460 181168 41472
rect 181088 41432 181168 41460
rect 181088 41404 181116 41432
rect 181162 41420 181168 41432
rect 181220 41420 181226 41472
rect 181070 41352 181076 41404
rect 181128 41352 181134 41404
rect 392670 41352 392676 41404
rect 392728 41392 392734 41404
rect 579890 41392 579896 41404
rect 392728 41364 579896 41392
rect 392728 41352 392734 41364
rect 579890 41352 579896 41364
rect 579948 41352 579954 41404
rect 219526 38740 219532 38752
rect 219487 38712 219532 38740
rect 219526 38700 219532 38712
rect 219584 38700 219590 38752
rect 239030 38740 239036 38752
rect 238991 38712 239036 38740
rect 239030 38700 239036 38712
rect 239088 38700 239094 38752
rect 168558 38632 168564 38684
rect 168616 38672 168622 38684
rect 168650 38672 168656 38684
rect 168616 38644 168656 38672
rect 168616 38632 168622 38644
rect 168650 38632 168656 38644
rect 168708 38632 168714 38684
rect 218238 38632 218244 38684
rect 218296 38672 218302 38684
rect 218330 38672 218336 38684
rect 218296 38644 218336 38672
rect 218296 38632 218302 38644
rect 218330 38632 218336 38644
rect 218388 38632 218394 38684
rect 256694 38632 256700 38684
rect 256752 38672 256758 38684
rect 256970 38672 256976 38684
rect 256752 38644 256976 38672
rect 256752 38632 256758 38644
rect 256970 38632 256976 38644
rect 257028 38632 257034 38684
rect 163130 38604 163136 38616
rect 163091 38576 163136 38604
rect 163130 38564 163136 38576
rect 163188 38564 163194 38616
rect 385313 38607 385371 38613
rect 385313 38573 385325 38607
rect 385359 38604 385371 38607
rect 385402 38604 385408 38616
rect 385359 38576 385408 38604
rect 385359 38573 385371 38576
rect 385313 38567 385371 38573
rect 385402 38564 385408 38576
rect 385460 38564 385466 38616
rect 182358 37312 182364 37324
rect 182319 37284 182364 37312
rect 182358 37272 182364 37284
rect 182416 37272 182422 37324
rect 210053 37315 210111 37321
rect 210053 37281 210065 37315
rect 210099 37312 210111 37315
rect 210142 37312 210148 37324
rect 210099 37284 210148 37312
rect 210099 37281 210111 37284
rect 210053 37275 210111 37281
rect 210142 37272 210148 37284
rect 210200 37272 210206 37324
rect 220998 37312 221004 37324
rect 220959 37284 221004 37312
rect 220998 37272 221004 37284
rect 221056 37272 221062 37324
rect 237282 37312 237288 37324
rect 237243 37284 237288 37312
rect 237282 37272 237288 37284
rect 237340 37272 237346 37324
rect 238662 37312 238668 37324
rect 238623 37284 238668 37312
rect 238662 37272 238668 37284
rect 238720 37272 238726 37324
rect 239030 37312 239036 37324
rect 238991 37284 239036 37312
rect 239030 37272 239036 37284
rect 239088 37272 239094 37324
rect 207382 37244 207388 37256
rect 207343 37216 207388 37244
rect 207382 37204 207388 37216
rect 207440 37204 207446 37256
rect 219526 35952 219532 35964
rect 219487 35924 219532 35952
rect 219526 35912 219532 35924
rect 219584 35912 219590 35964
rect 378134 35912 378140 35964
rect 378192 35952 378198 35964
rect 378318 35952 378324 35964
rect 378192 35924 378324 35952
rect 378192 35912 378198 35924
rect 378318 35912 378324 35924
rect 378376 35912 378382 35964
rect 3510 35844 3516 35896
rect 3568 35884 3574 35896
rect 152642 35884 152648 35896
rect 3568 35856 152648 35884
rect 3568 35844 3574 35856
rect 152642 35844 152648 35856
rect 152700 35844 152706 35896
rect 181070 34728 181076 34740
rect 181031 34700 181076 34728
rect 181070 34688 181076 34700
rect 181128 34688 181134 34740
rect 182358 31736 182364 31748
rect 182319 31708 182364 31736
rect 182358 31696 182364 31708
rect 182416 31696 182422 31748
rect 205726 31696 205732 31748
rect 205784 31736 205790 31748
rect 205910 31736 205916 31748
rect 205784 31708 205916 31736
rect 205784 31696 205790 31708
rect 205910 31696 205916 31708
rect 205968 31696 205974 31748
rect 225138 30336 225144 30388
rect 225196 30376 225202 30388
rect 225414 30376 225420 30388
rect 225196 30348 225420 30376
rect 225196 30336 225202 30348
rect 225414 30336 225420 30348
rect 225472 30336 225478 30388
rect 392578 30268 392584 30320
rect 392636 30308 392642 30320
rect 579890 30308 579896 30320
rect 392636 30280 579896 30308
rect 392636 30268 392642 30280
rect 579890 30268 579896 30280
rect 579948 30268 579954 30320
rect 159910 29588 159916 29640
rect 159968 29628 159974 29640
rect 218330 29628 218336 29640
rect 159968 29600 218336 29628
rect 159968 29588 159974 29600
rect 218330 29588 218336 29600
rect 218388 29588 218394 29640
rect 158898 29084 158904 29096
rect 158859 29056 158904 29084
rect 158898 29044 158904 29056
rect 158956 29044 158962 29096
rect 174262 29084 174268 29096
rect 174188 29056 174268 29084
rect 174188 29028 174216 29056
rect 174262 29044 174268 29056
rect 174320 29044 174326 29096
rect 163133 29019 163191 29025
rect 163133 28985 163145 29019
rect 163179 29016 163191 29019
rect 163222 29016 163228 29028
rect 163179 28988 163228 29016
rect 163179 28985 163191 28988
rect 163133 28979 163191 28985
rect 163222 28976 163228 28988
rect 163280 28976 163286 29028
rect 174170 28976 174176 29028
rect 174228 28976 174234 29028
rect 181073 29019 181131 29025
rect 181073 28985 181085 29019
rect 181119 29016 181131 29019
rect 181162 29016 181168 29028
rect 181119 28988 181168 29016
rect 181119 28985 181131 28988
rect 181073 28979 181131 28985
rect 181162 28976 181168 28988
rect 181220 28976 181226 29028
rect 182358 29016 182364 29028
rect 182319 28988 182364 29016
rect 182358 28976 182364 28988
rect 182416 28976 182422 29028
rect 216950 28976 216956 29028
rect 217008 29016 217014 29028
rect 217042 29016 217048 29028
rect 217008 28988 217048 29016
rect 217008 28976 217014 28988
rect 217042 28976 217048 28988
rect 217100 28976 217106 29028
rect 256510 28976 256516 29028
rect 256568 29016 256574 29028
rect 256786 29016 256792 29028
rect 256568 28988 256792 29016
rect 256568 28976 256574 28988
rect 256786 28976 256792 28988
rect 256844 28976 256850 29028
rect 385310 29016 385316 29028
rect 385271 28988 385316 29016
rect 385310 28976 385316 28988
rect 385368 28976 385374 29028
rect 222378 28908 222384 28960
rect 222436 28948 222442 28960
rect 222562 28948 222568 28960
rect 222436 28920 222568 28948
rect 222436 28908 222442 28920
rect 222562 28908 222568 28920
rect 222620 28908 222626 28960
rect 226610 28948 226616 28960
rect 226571 28920 226616 28948
rect 226610 28908 226616 28920
rect 226668 28908 226674 28960
rect 239030 28948 239036 28960
rect 238991 28920 239036 28948
rect 239030 28908 239036 28920
rect 239088 28908 239094 28960
rect 183462 28228 183468 28280
rect 183520 28268 183526 28280
rect 228082 28268 228088 28280
rect 183520 28240 228088 28268
rect 183520 28228 183526 28240
rect 228082 28228 228088 28240
rect 228140 28228 228146 28280
rect 183741 27727 183799 27733
rect 183741 27693 183753 27727
rect 183787 27724 183799 27727
rect 183922 27724 183928 27736
rect 183787 27696 183928 27724
rect 183787 27693 183799 27696
rect 183741 27687 183799 27693
rect 183922 27684 183928 27696
rect 183980 27684 183986 27736
rect 223942 27724 223948 27736
rect 223868 27696 223948 27724
rect 223868 27668 223896 27696
rect 223942 27684 223948 27696
rect 224000 27684 224006 27736
rect 207382 27656 207388 27668
rect 207343 27628 207388 27656
rect 207382 27616 207388 27628
rect 207440 27616 207446 27668
rect 223850 27616 223856 27668
rect 223908 27616 223914 27668
rect 158898 27588 158904 27600
rect 158859 27560 158904 27588
rect 158898 27548 158904 27560
rect 158956 27548 158962 27600
rect 181162 27588 181168 27600
rect 181123 27560 181168 27588
rect 181162 27548 181168 27560
rect 181220 27548 181226 27600
rect 216953 27591 217011 27597
rect 216953 27557 216965 27591
rect 216999 27588 217011 27591
rect 217042 27588 217048 27600
rect 216999 27560 217048 27588
rect 216999 27557 217011 27560
rect 216953 27551 217011 27557
rect 217042 27548 217048 27560
rect 217100 27548 217106 27600
rect 219526 27588 219532 27600
rect 219487 27560 219532 27588
rect 219526 27548 219532 27560
rect 219584 27548 219590 27600
rect 237282 27548 237288 27600
rect 237340 27548 237346 27600
rect 238662 27548 238668 27600
rect 238720 27548 238726 27600
rect 237193 27523 237251 27529
rect 237193 27489 237205 27523
rect 237239 27520 237251 27523
rect 237300 27520 237328 27548
rect 237239 27492 237328 27520
rect 238389 27523 238447 27529
rect 237239 27489 237251 27492
rect 237193 27483 237251 27489
rect 238389 27489 238401 27523
rect 238435 27520 238447 27523
rect 238680 27520 238708 27548
rect 238435 27492 238708 27520
rect 238435 27489 238447 27492
rect 238389 27483 238447 27489
rect 186222 26868 186228 26920
rect 186280 26908 186286 26920
rect 229278 26908 229284 26920
rect 186280 26880 229284 26908
rect 186280 26868 186286 26880
rect 229278 26868 229284 26880
rect 229336 26868 229342 26920
rect 183738 26364 183744 26376
rect 183699 26336 183744 26364
rect 183738 26324 183744 26336
rect 183796 26324 183802 26376
rect 183738 26228 183744 26240
rect 183699 26200 183744 26228
rect 183738 26188 183744 26200
rect 183796 26188 183802 26240
rect 157242 25508 157248 25560
rect 157300 25548 157306 25560
rect 215938 25548 215944 25560
rect 157300 25520 215944 25548
rect 157300 25508 157306 25520
rect 215938 25508 215944 25520
rect 215996 25508 216002 25560
rect 153102 24080 153108 24132
rect 153160 24120 153166 24132
rect 214558 24120 214564 24132
rect 153160 24092 214564 24120
rect 153160 24080 153166 24092
rect 214558 24080 214564 24092
rect 214616 24080 214622 24132
rect 141970 22720 141976 22772
rect 142028 22760 142034 22772
rect 211246 22760 211252 22772
rect 142028 22732 211252 22760
rect 142028 22720 142034 22732
rect 211246 22720 211252 22732
rect 211304 22720 211310 22772
rect 239030 22760 239036 22772
rect 238991 22732 239036 22760
rect 239030 22720 239036 22732
rect 239088 22720 239094 22772
rect 182358 22108 182364 22160
rect 182416 22108 182422 22160
rect 207201 22151 207259 22157
rect 207201 22117 207213 22151
rect 207247 22148 207259 22151
rect 207382 22148 207388 22160
rect 207247 22120 207388 22148
rect 207247 22117 207259 22120
rect 207201 22111 207259 22117
rect 207382 22108 207388 22120
rect 207440 22108 207446 22160
rect 221090 22108 221096 22160
rect 221148 22108 221154 22160
rect 156230 22040 156236 22092
rect 156288 22080 156294 22092
rect 156414 22080 156420 22092
rect 156288 22052 156420 22080
rect 156288 22040 156294 22052
rect 156414 22040 156420 22052
rect 156472 22040 156478 22092
rect 182376 22012 182404 22108
rect 200298 22040 200304 22092
rect 200356 22040 200362 22092
rect 182450 22012 182456 22024
rect 182376 21984 182456 22012
rect 182450 21972 182456 21984
rect 182508 21972 182514 22024
rect 200316 22012 200344 22040
rect 221108 22024 221136 22108
rect 256878 22040 256884 22092
rect 256936 22080 256942 22092
rect 257062 22080 257068 22092
rect 256936 22052 257068 22080
rect 256936 22040 256942 22052
rect 257062 22040 257068 22052
rect 257120 22040 257126 22092
rect 200390 22012 200396 22024
rect 200316 21984 200396 22012
rect 200390 21972 200396 21984
rect 200448 21972 200454 22024
rect 221090 21972 221096 22024
rect 221148 21972 221154 22024
rect 188982 21360 188988 21412
rect 189040 21400 189046 21412
rect 230658 21400 230664 21412
rect 189040 21372 230664 21400
rect 189040 21360 189046 21372
rect 230658 21360 230664 21372
rect 230716 21360 230722 21412
rect 292298 21360 292304 21412
rect 292356 21400 292362 21412
rect 339586 21400 339592 21412
rect 292356 21372 339592 21400
rect 292356 21360 292362 21372
rect 339586 21360 339592 21372
rect 339644 21360 339650 21412
rect 365530 21360 365536 21412
rect 365588 21400 365594 21412
rect 520366 21400 520372 21412
rect 365588 21372 520372 21400
rect 365588 21360 365594 21372
rect 520366 21360 520372 21372
rect 520424 21360 520430 21412
rect 180702 19932 180708 19984
rect 180760 19972 180766 19984
rect 226613 19975 226671 19981
rect 226613 19972 226625 19975
rect 180760 19944 226625 19972
rect 180760 19932 180766 19944
rect 226613 19941 226625 19944
rect 226659 19941 226671 19975
rect 226613 19935 226671 19941
rect 291010 19932 291016 19984
rect 291068 19972 291074 19984
rect 336734 19972 336740 19984
rect 291068 19944 336740 19972
rect 291068 19932 291074 19944
rect 336734 19932 336740 19944
rect 336792 19932 336798 19984
rect 361482 19932 361488 19984
rect 361540 19972 361546 19984
rect 510614 19972 510620 19984
rect 361540 19944 510620 19972
rect 361540 19932 361546 19944
rect 510614 19932 510620 19944
rect 510672 19932 510678 19984
rect 156414 19292 156420 19304
rect 156375 19264 156420 19292
rect 156414 19252 156420 19264
rect 156472 19252 156478 19304
rect 200390 19292 200396 19304
rect 200351 19264 200396 19292
rect 200390 19252 200396 19264
rect 200448 19252 200454 19304
rect 222470 19292 222476 19304
rect 222431 19264 222476 19292
rect 222470 19252 222476 19264
rect 222528 19252 222534 19304
rect 257062 19292 257068 19304
rect 257023 19264 257068 19292
rect 257062 19252 257068 19264
rect 257120 19252 257126 19304
rect 385037 19295 385095 19301
rect 385037 19261 385049 19295
rect 385083 19292 385095 19295
rect 385126 19292 385132 19304
rect 385083 19264 385132 19292
rect 385083 19261 385095 19264
rect 385037 19255 385095 19261
rect 385126 19252 385132 19264
rect 385184 19252 385190 19304
rect 158898 19224 158904 19236
rect 158859 19196 158904 19224
rect 158898 19184 158904 19196
rect 158956 19184 158962 19236
rect 173802 18572 173808 18624
rect 173860 18612 173866 18624
rect 223850 18612 223856 18624
rect 173860 18584 223856 18612
rect 173860 18572 173866 18584
rect 223850 18572 223856 18584
rect 223908 18572 223914 18624
rect 286778 18572 286784 18624
rect 286836 18612 286842 18624
rect 325694 18612 325700 18624
rect 286836 18584 325700 18612
rect 286836 18572 286842 18584
rect 325694 18572 325700 18584
rect 325752 18572 325758 18624
rect 360102 18572 360108 18624
rect 360160 18612 360166 18624
rect 506474 18612 506480 18624
rect 360160 18584 506480 18612
rect 360160 18572 360166 18584
rect 506474 18572 506480 18584
rect 506532 18572 506538 18624
rect 181162 18000 181168 18012
rect 181123 17972 181168 18000
rect 181162 17960 181168 17972
rect 181220 17960 181226 18012
rect 185118 17960 185124 18012
rect 185176 18000 185182 18012
rect 185394 18000 185400 18012
rect 185176 17972 185400 18000
rect 185176 17960 185182 17972
rect 185394 17960 185400 17972
rect 185452 17960 185458 18012
rect 207198 18000 207204 18012
rect 207159 17972 207204 18000
rect 207198 17960 207204 17972
rect 207256 17960 207262 18012
rect 135162 17212 135168 17264
rect 135220 17252 135226 17264
rect 208394 17252 208400 17264
rect 135220 17224 208400 17252
rect 135220 17212 135226 17224
rect 208394 17212 208400 17224
rect 208452 17212 208458 17264
rect 281350 17212 281356 17264
rect 281408 17252 281414 17264
rect 311894 17252 311900 17264
rect 281408 17224 311900 17252
rect 281408 17212 281414 17224
rect 311894 17212 311900 17224
rect 311952 17212 311958 17264
rect 358722 17212 358728 17264
rect 358780 17252 358786 17264
rect 502426 17252 502432 17264
rect 358780 17224 502432 17252
rect 358780 17212 358786 17224
rect 502426 17212 502432 17224
rect 502484 17212 502490 17264
rect 183738 16640 183744 16652
rect 183699 16612 183744 16640
rect 183738 16600 183744 16612
rect 183796 16600 183802 16652
rect 378134 16600 378140 16652
rect 378192 16640 378198 16652
rect 378318 16640 378324 16652
rect 378192 16612 378324 16640
rect 378192 16600 378198 16612
rect 378318 16600 378324 16612
rect 378376 16600 378382 16652
rect 187602 15852 187608 15904
rect 187660 15892 187666 15904
rect 229186 15892 229192 15904
rect 187660 15864 229192 15892
rect 187660 15852 187666 15864
rect 229186 15852 229192 15864
rect 229244 15852 229250 15904
rect 277118 15852 277124 15904
rect 277176 15892 277182 15904
rect 300854 15892 300860 15904
rect 277176 15864 300860 15892
rect 277176 15852 277182 15864
rect 300854 15852 300860 15864
rect 300912 15852 300918 15904
rect 357342 15852 357348 15904
rect 357400 15892 357406 15904
rect 499574 15892 499580 15904
rect 357400 15864 499580 15892
rect 357400 15852 357406 15864
rect 499574 15852 499580 15864
rect 499632 15852 499638 15904
rect 180978 14492 180984 14544
rect 181036 14532 181042 14544
rect 181162 14532 181168 14544
rect 181036 14504 181168 14532
rect 181036 14492 181042 14504
rect 181162 14492 181168 14504
rect 181220 14492 181226 14544
rect 184842 14424 184848 14476
rect 184900 14464 184906 14476
rect 227806 14464 227812 14476
rect 184900 14436 227812 14464
rect 184900 14424 184906 14436
rect 227806 14424 227812 14436
rect 227864 14424 227870 14476
rect 285398 14424 285404 14476
rect 285456 14464 285462 14476
rect 321646 14464 321652 14476
rect 285456 14436 321652 14464
rect 285456 14424 285462 14436
rect 321646 14424 321652 14436
rect 321704 14424 321710 14476
rect 354582 14424 354588 14476
rect 354640 14464 354646 14476
rect 494146 14464 494152 14476
rect 354640 14436 494152 14464
rect 354640 14424 354646 14436
rect 494146 14424 494152 14436
rect 494204 14424 494210 14476
rect 183738 13172 183744 13184
rect 183699 13144 183744 13172
rect 183738 13132 183744 13144
rect 183796 13132 183802 13184
rect 278590 13132 278596 13184
rect 278648 13172 278654 13184
rect 304994 13172 305000 13184
rect 278648 13144 305000 13172
rect 278648 13132 278654 13144
rect 304994 13132 305000 13144
rect 305052 13132 305058 13184
rect 176562 13064 176568 13116
rect 176620 13104 176626 13116
rect 225138 13104 225144 13116
rect 176620 13076 225144 13104
rect 176620 13064 176626 13076
rect 225138 13064 225144 13076
rect 225196 13064 225202 13116
rect 282638 13064 282644 13116
rect 282696 13104 282702 13116
rect 314654 13104 314660 13116
rect 282696 13076 314660 13104
rect 282696 13064 282702 13076
rect 314654 13064 314660 13076
rect 314712 13064 314718 13116
rect 355962 13064 355968 13116
rect 356020 13104 356026 13116
rect 495434 13104 495440 13116
rect 356020 13076 495440 13104
rect 356020 13064 356026 13076
rect 495434 13064 495440 13076
rect 495492 13064 495498 13116
rect 185118 12492 185124 12504
rect 185079 12464 185124 12492
rect 185118 12452 185124 12464
rect 185176 12452 185182 12504
rect 156414 12424 156420 12436
rect 156375 12396 156420 12424
rect 156414 12384 156420 12396
rect 156472 12384 156478 12436
rect 205726 12384 205732 12436
rect 205784 12424 205790 12436
rect 205910 12424 205916 12436
rect 205784 12396 205916 12424
rect 205784 12384 205790 12396
rect 205910 12384 205916 12396
rect 205968 12384 205974 12436
rect 257062 12288 257068 12300
rect 257023 12260 257068 12288
rect 257062 12248 257068 12260
rect 257120 12248 257126 12300
rect 279970 11772 279976 11824
rect 280028 11812 280034 11824
rect 307754 11812 307760 11824
rect 280028 11784 307760 11812
rect 280028 11772 280034 11784
rect 307754 11772 307760 11784
rect 307812 11772 307818 11824
rect 23382 11704 23388 11756
rect 23440 11744 23446 11756
rect 164326 11744 164332 11756
rect 23440 11716 164332 11744
rect 23440 11704 23446 11716
rect 164326 11704 164332 11716
rect 164384 11704 164390 11756
rect 169386 11704 169392 11756
rect 169444 11744 169450 11756
rect 222473 11747 222531 11753
rect 222473 11744 222485 11747
rect 169444 11716 222485 11744
rect 169444 11704 169450 11716
rect 222473 11713 222485 11716
rect 222519 11713 222531 11747
rect 222473 11707 222531 11713
rect 289538 11704 289544 11756
rect 289596 11744 289602 11756
rect 332594 11744 332600 11756
rect 289596 11716 332600 11744
rect 289596 11704 289602 11716
rect 332594 11704 332600 11716
rect 332652 11704 332658 11756
rect 351730 11704 351736 11756
rect 351788 11744 351794 11756
rect 485866 11744 485872 11756
rect 351788 11716 485872 11744
rect 351788 11704 351794 11716
rect 485866 11704 485872 11716
rect 485924 11704 485930 11756
rect 192018 10344 192024 10396
rect 192076 10384 192082 10396
rect 231946 10384 231952 10396
rect 192076 10356 231952 10384
rect 192076 10344 192082 10356
rect 231946 10344 231952 10356
rect 232004 10344 232010 10396
rect 278682 10344 278688 10396
rect 278740 10384 278746 10396
rect 305086 10384 305092 10396
rect 278740 10356 305092 10384
rect 278740 10344 278746 10356
rect 305086 10344 305092 10356
rect 305144 10344 305150 10396
rect 13630 10276 13636 10328
rect 13688 10316 13694 10328
rect 160186 10316 160192 10328
rect 13688 10288 160192 10316
rect 13688 10276 13694 10288
rect 160186 10276 160192 10288
rect 160244 10276 160250 10328
rect 165890 10276 165896 10328
rect 165948 10316 165954 10328
rect 221090 10316 221096 10328
rect 165948 10288 221096 10316
rect 165948 10276 165954 10288
rect 221090 10276 221096 10288
rect 221148 10276 221154 10328
rect 288250 10276 288256 10328
rect 288308 10316 288314 10328
rect 329834 10316 329840 10328
rect 288308 10288 329840 10316
rect 288308 10276 288314 10288
rect 329834 10276 329840 10288
rect 329892 10276 329898 10328
rect 353202 10276 353208 10328
rect 353260 10316 353266 10328
rect 488534 10316 488540 10328
rect 353260 10288 488540 10316
rect 353260 10276 353266 10288
rect 488534 10276 488540 10288
rect 488592 10276 488598 10328
rect 158898 9664 158904 9716
rect 158956 9704 158962 9716
rect 158990 9704 158996 9716
rect 158956 9676 158996 9704
rect 158956 9664 158962 9676
rect 158990 9664 158996 9676
rect 159048 9664 159054 9716
rect 200390 9704 200396 9716
rect 200351 9676 200396 9704
rect 200390 9664 200396 9676
rect 200448 9664 200454 9716
rect 216950 9704 216956 9716
rect 216911 9676 216956 9704
rect 216950 9664 216956 9676
rect 217008 9664 217014 9716
rect 219526 9704 219532 9716
rect 219487 9676 219532 9704
rect 219526 9664 219532 9676
rect 219584 9664 219590 9716
rect 237190 9704 237196 9716
rect 237151 9676 237196 9704
rect 237190 9664 237196 9676
rect 237248 9664 237254 9716
rect 238386 9704 238392 9716
rect 238347 9676 238392 9704
rect 238386 9664 238392 9676
rect 238444 9664 238450 9716
rect 385034 9704 385040 9716
rect 384995 9676 385040 9704
rect 385034 9664 385040 9676
rect 385092 9664 385098 9716
rect 312538 9596 312544 9648
rect 312596 9636 312602 9648
rect 313366 9636 313372 9648
rect 312596 9608 313372 9636
rect 312596 9596 312602 9608
rect 313366 9596 313372 9608
rect 313424 9596 313430 9648
rect 326890 9596 326896 9648
rect 326948 9636 326954 9648
rect 423950 9636 423956 9648
rect 326948 9608 423956 9636
rect 326948 9596 326954 9608
rect 423950 9596 423956 9608
rect 424008 9596 424014 9648
rect 328178 9528 328184 9580
rect 328236 9568 328242 9580
rect 427538 9568 427544 9580
rect 328236 9540 427544 9568
rect 328236 9528 328242 9540
rect 427538 9528 427544 9540
rect 427596 9528 427602 9580
rect 329650 9460 329656 9512
rect 329708 9500 329714 9512
rect 431126 9500 431132 9512
rect 329708 9472 431132 9500
rect 329708 9460 329714 9472
rect 431126 9460 431132 9472
rect 431184 9460 431190 9512
rect 330938 9392 330944 9444
rect 330996 9432 331002 9444
rect 434622 9432 434628 9444
rect 330996 9404 434628 9432
rect 330996 9392 331002 9404
rect 434622 9392 434628 9404
rect 434680 9392 434686 9444
rect 332410 9324 332416 9376
rect 332468 9364 332474 9376
rect 438210 9364 438216 9376
rect 332468 9336 438216 9364
rect 332468 9324 332474 9336
rect 438210 9324 438216 9336
rect 438268 9324 438274 9376
rect 333698 9256 333704 9308
rect 333756 9296 333762 9308
rect 441798 9296 441804 9308
rect 333756 9268 441804 9296
rect 333756 9256 333762 9268
rect 441798 9256 441804 9268
rect 441856 9256 441862 9308
rect 335170 9188 335176 9240
rect 335228 9228 335234 9240
rect 445386 9228 445392 9240
rect 335228 9200 445392 9228
rect 335228 9188 335234 9200
rect 445386 9188 445392 9200
rect 445444 9188 445450 9240
rect 336550 9120 336556 9172
rect 336608 9160 336614 9172
rect 448974 9160 448980 9172
rect 336608 9132 448980 9160
rect 336608 9120 336614 9132
rect 448974 9120 448980 9132
rect 449032 9120 449038 9172
rect 337930 9052 337936 9104
rect 337988 9092 337994 9104
rect 452470 9092 452476 9104
rect 337988 9064 452476 9092
rect 337988 9052 337994 9064
rect 452470 9052 452476 9064
rect 452528 9052 452534 9104
rect 184750 8984 184756 9036
rect 184808 9024 184814 9036
rect 229094 9024 229100 9036
rect 184808 8996 229100 9024
rect 184808 8984 184814 8996
rect 229094 8984 229100 8996
rect 229152 8984 229158 9036
rect 278038 8984 278044 9036
rect 278096 9024 278102 9036
rect 299106 9024 299112 9036
rect 278096 8996 299112 9024
rect 278096 8984 278102 8996
rect 299106 8984 299112 8996
rect 299164 8984 299170 9036
rect 339218 8984 339224 9036
rect 339276 9024 339282 9036
rect 456058 9024 456064 9036
rect 339276 8996 456064 9024
rect 339276 8984 339282 8996
rect 456058 8984 456064 8996
rect 456116 8984 456122 9036
rect 162302 8916 162308 8968
rect 162360 8956 162366 8968
rect 219526 8956 219532 8968
rect 162360 8928 219532 8956
rect 162360 8916 162366 8928
rect 219526 8916 219532 8928
rect 219584 8916 219590 8968
rect 275830 8916 275836 8968
rect 275888 8956 275894 8968
rect 297726 8956 297732 8968
rect 275888 8928 297732 8956
rect 275888 8916 275894 8928
rect 297726 8916 297732 8928
rect 297784 8916 297790 8968
rect 340690 8916 340696 8968
rect 340748 8956 340754 8968
rect 459646 8956 459652 8968
rect 340748 8928 459652 8956
rect 340748 8916 340754 8928
rect 459646 8916 459652 8928
rect 459704 8916 459710 8968
rect 324222 8848 324228 8900
rect 324280 8888 324286 8900
rect 420362 8888 420368 8900
rect 324280 8860 420368 8888
rect 324280 8848 324286 8860
rect 420362 8848 420368 8860
rect 420420 8848 420426 8900
rect 322750 8780 322756 8832
rect 322808 8820 322814 8832
rect 416866 8820 416872 8832
rect 322808 8792 416872 8820
rect 322808 8780 322814 8792
rect 416866 8780 416872 8792
rect 416924 8780 416930 8832
rect 321462 8712 321468 8764
rect 321520 8752 321526 8764
rect 413278 8752 413284 8764
rect 321520 8724 413284 8752
rect 321520 8712 321526 8724
rect 413278 8712 413284 8724
rect 413336 8712 413342 8764
rect 319990 8644 319996 8696
rect 320048 8684 320054 8696
rect 409690 8684 409696 8696
rect 320048 8656 409696 8684
rect 320048 8644 320054 8656
rect 409690 8644 409696 8656
rect 409748 8644 409754 8696
rect 318702 8576 318708 8628
rect 318760 8616 318766 8628
rect 406102 8616 406108 8628
rect 318760 8588 406108 8616
rect 318760 8576 318766 8588
rect 406102 8576 406108 8588
rect 406160 8576 406166 8628
rect 317230 8508 317236 8560
rect 317288 8548 317294 8560
rect 402514 8548 402520 8560
rect 317288 8520 402520 8548
rect 317288 8508 317294 8520
rect 402514 8508 402520 8520
rect 402572 8508 402578 8560
rect 315942 8440 315948 8492
rect 316000 8480 316006 8492
rect 399018 8480 399024 8492
rect 316000 8452 399024 8480
rect 316000 8440 316006 8452
rect 399018 8440 399024 8452
rect 399076 8440 399082 8492
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 152458 8276 152464 8288
rect 3476 8248 152464 8276
rect 3476 8236 3482 8248
rect 152458 8236 152464 8248
rect 152516 8236 152522 8288
rect 375098 8236 375104 8288
rect 375156 8276 375162 8288
rect 545298 8276 545304 8288
rect 375156 8248 545304 8276
rect 375156 8236 375162 8248
rect 545298 8236 545304 8248
rect 545356 8236 545362 8288
rect 94498 8168 94504 8220
rect 94556 8208 94562 8220
rect 191926 8208 191932 8220
rect 94556 8180 191932 8208
rect 94556 8168 94562 8180
rect 191926 8168 191932 8180
rect 191984 8168 191990 8220
rect 299198 8168 299204 8220
rect 299256 8208 299262 8220
rect 356146 8208 356152 8220
rect 299256 8180 356152 8208
rect 299256 8168 299262 8180
rect 356146 8168 356152 8180
rect 356204 8168 356210 8220
rect 376478 8168 376484 8220
rect 376536 8208 376542 8220
rect 548886 8208 548892 8220
rect 376536 8180 548892 8208
rect 376536 8168 376542 8180
rect 548886 8168 548892 8180
rect 548944 8168 548950 8220
rect 77846 8100 77852 8152
rect 77904 8140 77910 8152
rect 186498 8140 186504 8152
rect 77904 8112 186504 8140
rect 77904 8100 77910 8112
rect 186498 8100 186504 8112
rect 186556 8100 186562 8152
rect 300578 8100 300584 8152
rect 300636 8140 300642 8152
rect 359734 8140 359740 8152
rect 300636 8112 359740 8140
rect 300636 8100 300642 8112
rect 359734 8100 359740 8112
rect 359792 8100 359798 8152
rect 377858 8100 377864 8152
rect 377916 8140 377922 8152
rect 552382 8140 552388 8152
rect 377916 8112 552388 8140
rect 377916 8100 377922 8112
rect 552382 8100 552388 8112
rect 552440 8100 552446 8152
rect 74258 8032 74264 8084
rect 74316 8072 74322 8084
rect 183741 8075 183799 8081
rect 183741 8072 183753 8075
rect 74316 8044 183753 8072
rect 74316 8032 74322 8044
rect 183741 8041 183753 8044
rect 183787 8041 183799 8075
rect 183741 8035 183799 8041
rect 302050 8032 302056 8084
rect 302108 8072 302114 8084
rect 363322 8072 363328 8084
rect 302108 8044 363328 8072
rect 302108 8032 302114 8044
rect 363322 8032 363328 8044
rect 363380 8032 363386 8084
rect 379238 8032 379244 8084
rect 379296 8072 379302 8084
rect 555970 8072 555976 8084
rect 379296 8044 555976 8072
rect 379296 8032 379302 8044
rect 555970 8032 555976 8044
rect 556028 8032 556034 8084
rect 70670 7964 70676 8016
rect 70728 8004 70734 8016
rect 182358 8004 182364 8016
rect 70728 7976 182364 8004
rect 70728 7964 70734 7976
rect 182358 7964 182364 7976
rect 182416 7964 182422 8016
rect 303338 7964 303344 8016
rect 303396 8004 303402 8016
rect 366910 8004 366916 8016
rect 303396 7976 366916 8004
rect 303396 7964 303402 7976
rect 366910 7964 366916 7976
rect 366968 7964 366974 8016
rect 380618 7964 380624 8016
rect 380676 8004 380682 8016
rect 559558 8004 559564 8016
rect 380676 7976 559564 8004
rect 380676 7964 380682 7976
rect 559558 7964 559564 7976
rect 559616 7964 559622 8016
rect 67174 7896 67180 7948
rect 67232 7936 67238 7948
rect 180978 7936 180984 7948
rect 67232 7908 180984 7936
rect 67232 7896 67238 7908
rect 180978 7896 180984 7908
rect 181036 7896 181042 7948
rect 304718 7896 304724 7948
rect 304776 7936 304782 7948
rect 370406 7936 370412 7948
rect 304776 7908 370412 7936
rect 304776 7896 304782 7908
rect 370406 7896 370412 7908
rect 370464 7896 370470 7948
rect 381998 7896 382004 7948
rect 382056 7936 382062 7948
rect 563146 7936 563152 7948
rect 382056 7908 563152 7936
rect 382056 7896 382062 7908
rect 563146 7896 563152 7908
rect 563204 7896 563210 7948
rect 63586 7828 63592 7880
rect 63644 7868 63650 7880
rect 179506 7868 179512 7880
rect 63644 7840 179512 7868
rect 63644 7828 63650 7840
rect 179506 7828 179512 7840
rect 179564 7828 179570 7880
rect 306098 7828 306104 7880
rect 306156 7868 306162 7880
rect 373994 7868 374000 7880
rect 306156 7840 374000 7868
rect 306156 7828 306162 7840
rect 373994 7828 374000 7840
rect 374052 7828 374058 7880
rect 383470 7828 383476 7880
rect 383528 7868 383534 7880
rect 566734 7868 566740 7880
rect 383528 7840 566740 7868
rect 383528 7828 383534 7840
rect 566734 7828 566740 7840
rect 566792 7828 566798 7880
rect 59998 7760 60004 7812
rect 60056 7800 60062 7812
rect 178126 7800 178132 7812
rect 60056 7772 178132 7800
rect 60056 7760 60062 7772
rect 178126 7760 178132 7772
rect 178184 7760 178190 7812
rect 307570 7760 307576 7812
rect 307628 7800 307634 7812
rect 377582 7800 377588 7812
rect 307628 7772 377588 7800
rect 307628 7760 307634 7772
rect 377582 7760 377588 7772
rect 377640 7760 377646 7812
rect 384758 7760 384764 7812
rect 384816 7800 384822 7812
rect 570230 7800 570236 7812
rect 384816 7772 570236 7800
rect 384816 7760 384822 7772
rect 570230 7760 570236 7772
rect 570288 7760 570294 7812
rect 56410 7692 56416 7744
rect 56468 7732 56474 7744
rect 176746 7732 176752 7744
rect 56468 7704 176752 7732
rect 56468 7692 56474 7704
rect 176746 7692 176752 7704
rect 176804 7692 176810 7744
rect 308858 7692 308864 7744
rect 308916 7732 308922 7744
rect 381170 7732 381176 7744
rect 308916 7704 381176 7732
rect 308916 7692 308922 7704
rect 381170 7692 381176 7704
rect 381228 7692 381234 7744
rect 386138 7692 386144 7744
rect 386196 7732 386202 7744
rect 573818 7732 573824 7744
rect 386196 7704 573824 7732
rect 386196 7692 386202 7704
rect 573818 7692 573824 7704
rect 573876 7692 573882 7744
rect 52822 7624 52828 7676
rect 52880 7664 52886 7676
rect 175366 7664 175372 7676
rect 52880 7636 175372 7664
rect 52880 7624 52886 7636
rect 175366 7624 175372 7636
rect 175424 7624 175430 7676
rect 271598 7624 271604 7676
rect 271656 7664 271662 7676
rect 287146 7664 287152 7676
rect 271656 7636 287152 7664
rect 271656 7624 271662 7636
rect 287146 7624 287152 7636
rect 287204 7624 287210 7676
rect 310330 7624 310336 7676
rect 310388 7664 310394 7676
rect 384666 7664 384672 7676
rect 310388 7636 384672 7664
rect 310388 7624 310394 7636
rect 384666 7624 384672 7636
rect 384724 7624 384730 7676
rect 387518 7624 387524 7676
rect 387576 7664 387582 7676
rect 577406 7664 577412 7676
rect 387576 7636 577412 7664
rect 387576 7624 387582 7636
rect 577406 7624 577412 7636
rect 577464 7624 577470 7676
rect 49326 7556 49332 7608
rect 49384 7596 49390 7608
rect 174078 7596 174084 7608
rect 49384 7568 174084 7596
rect 49384 7556 49390 7568
rect 174078 7556 174084 7568
rect 174136 7556 174142 7608
rect 201494 7556 201500 7608
rect 201552 7596 201558 7608
rect 236086 7596 236092 7608
rect 201552 7568 236092 7596
rect 201552 7556 201558 7568
rect 236086 7556 236092 7568
rect 236144 7556 236150 7608
rect 274450 7556 274456 7608
rect 274508 7596 274514 7608
rect 295518 7596 295524 7608
rect 274508 7568 295524 7596
rect 274508 7556 274514 7568
rect 295518 7556 295524 7568
rect 295576 7556 295582 7608
rect 311618 7556 311624 7608
rect 311676 7596 311682 7608
rect 388254 7596 388260 7608
rect 311676 7568 388260 7596
rect 311676 7556 311682 7568
rect 388254 7556 388260 7568
rect 388312 7556 388318 7608
rect 388898 7556 388904 7608
rect 388956 7596 388962 7608
rect 580994 7596 581000 7608
rect 388956 7568 581000 7596
rect 388956 7556 388962 7568
rect 580994 7556 581000 7568
rect 581052 7556 581058 7608
rect 98086 7488 98092 7540
rect 98144 7528 98150 7540
rect 193306 7528 193312 7540
rect 98144 7500 193312 7528
rect 98144 7488 98150 7500
rect 193306 7488 193312 7500
rect 193364 7488 193370 7540
rect 373810 7488 373816 7540
rect 373868 7528 373874 7540
rect 541710 7528 541716 7540
rect 373868 7500 541716 7528
rect 373868 7488 373874 7500
rect 541710 7488 541716 7500
rect 541768 7488 541774 7540
rect 101582 7420 101588 7472
rect 101640 7460 101646 7472
rect 194686 7460 194692 7472
rect 101640 7432 194692 7460
rect 101640 7420 101646 7432
rect 194686 7420 194692 7432
rect 194744 7420 194750 7472
rect 372522 7420 372528 7472
rect 372580 7460 372586 7472
rect 538122 7460 538128 7472
rect 372580 7432 538128 7460
rect 372580 7420 372586 7432
rect 538122 7420 538128 7432
rect 538180 7420 538186 7472
rect 105170 7352 105176 7404
rect 105228 7392 105234 7404
rect 197446 7392 197452 7404
rect 105228 7364 197452 7392
rect 105228 7352 105234 7364
rect 197446 7352 197452 7364
rect 197504 7352 197510 7404
rect 371050 7352 371056 7404
rect 371108 7392 371114 7404
rect 534534 7392 534540 7404
rect 371108 7364 534540 7392
rect 371108 7352 371114 7364
rect 534534 7352 534540 7364
rect 534592 7352 534598 7404
rect 108758 7284 108764 7336
rect 108816 7324 108822 7336
rect 198918 7324 198924 7336
rect 108816 7296 198924 7324
rect 108816 7284 108822 7296
rect 198918 7284 198924 7296
rect 198976 7284 198982 7336
rect 369670 7284 369676 7336
rect 369728 7324 369734 7336
rect 531038 7324 531044 7336
rect 369728 7296 531044 7324
rect 369728 7284 369734 7296
rect 531038 7284 531044 7296
rect 531096 7284 531102 7336
rect 112346 7216 112352 7268
rect 112404 7256 112410 7268
rect 200206 7256 200212 7268
rect 112404 7228 200212 7256
rect 112404 7216 112410 7228
rect 200206 7216 200212 7228
rect 200264 7216 200270 7268
rect 368290 7216 368296 7268
rect 368348 7256 368354 7268
rect 527450 7256 527456 7268
rect 368348 7228 527456 7256
rect 368348 7216 368354 7228
rect 527450 7216 527456 7228
rect 527508 7216 527514 7268
rect 115934 7148 115940 7200
rect 115992 7188 115998 7200
rect 201678 7188 201684 7200
rect 115992 7160 201684 7188
rect 115992 7148 115998 7160
rect 201678 7148 201684 7160
rect 201736 7148 201742 7200
rect 366818 7148 366824 7200
rect 366876 7188 366882 7200
rect 523862 7188 523868 7200
rect 366876 7160 523868 7188
rect 366876 7148 366882 7160
rect 523862 7148 523868 7160
rect 523920 7148 523926 7200
rect 119430 7080 119436 7132
rect 119488 7120 119494 7132
rect 203058 7120 203064 7132
rect 119488 7092 203064 7120
rect 119488 7080 119494 7092
rect 203058 7080 203064 7092
rect 203116 7080 203122 7132
rect 314470 7080 314476 7132
rect 314528 7120 314534 7132
rect 395430 7120 395436 7132
rect 314528 7092 395436 7120
rect 314528 7080 314534 7092
rect 395430 7080 395436 7092
rect 395488 7080 395494 7132
rect 123018 7012 123024 7064
rect 123076 7052 123082 7064
rect 204346 7052 204352 7064
rect 123076 7024 204352 7052
rect 123076 7012 123082 7024
rect 204346 7012 204352 7024
rect 204404 7012 204410 7064
rect 313182 7012 313188 7064
rect 313240 7052 313246 7064
rect 391842 7052 391848 7064
rect 313240 7024 391848 7052
rect 313240 7012 313246 7024
rect 391842 7012 391848 7024
rect 391900 7012 391906 7064
rect 132586 6808 132592 6860
rect 132644 6848 132650 6860
rect 207290 6848 207296 6860
rect 132644 6820 207296 6848
rect 132644 6808 132650 6820
rect 207290 6808 207296 6820
rect 207348 6808 207354 6860
rect 338022 6808 338028 6860
rect 338080 6848 338086 6860
rect 451274 6848 451280 6860
rect 338080 6820 451280 6848
rect 338080 6808 338086 6820
rect 451274 6808 451280 6820
rect 451332 6808 451338 6860
rect 128998 6740 129004 6792
rect 129056 6780 129062 6792
rect 205726 6780 205732 6792
rect 129056 6752 205732 6780
rect 129056 6740 129062 6752
rect 205726 6740 205732 6752
rect 205784 6740 205790 6792
rect 339310 6740 339316 6792
rect 339368 6780 339374 6792
rect 454862 6780 454868 6792
rect 339368 6752 454868 6780
rect 339368 6740 339374 6752
rect 454862 6740 454868 6752
rect 454920 6740 454926 6792
rect 90910 6672 90916 6724
rect 90968 6712 90974 6724
rect 190546 6712 190552 6724
rect 90968 6684 190552 6712
rect 90968 6672 90974 6684
rect 190546 6672 190552 6684
rect 190604 6672 190610 6724
rect 340782 6672 340788 6724
rect 340840 6712 340846 6724
rect 458450 6712 458456 6724
rect 340840 6684 458456 6712
rect 340840 6672 340846 6684
rect 458450 6672 458456 6684
rect 458508 6672 458514 6724
rect 87322 6604 87328 6656
rect 87380 6644 87386 6656
rect 189166 6644 189172 6656
rect 87380 6616 189172 6644
rect 87380 6604 87386 6616
rect 189166 6604 189172 6616
rect 189224 6604 189230 6656
rect 342070 6604 342076 6656
rect 342128 6644 342134 6656
rect 462038 6644 462044 6656
rect 342128 6616 462044 6644
rect 342128 6604 342134 6616
rect 462038 6604 462044 6616
rect 462096 6604 462102 6656
rect 83826 6536 83832 6588
rect 83884 6576 83890 6588
rect 187786 6576 187792 6588
rect 83884 6548 187792 6576
rect 83884 6536 83890 6548
rect 187786 6536 187792 6548
rect 187844 6536 187850 6588
rect 343542 6536 343548 6588
rect 343600 6576 343606 6588
rect 465626 6576 465632 6588
rect 343600 6548 465632 6576
rect 343600 6536 343606 6548
rect 465626 6536 465632 6548
rect 465684 6536 465690 6588
rect 44542 6468 44548 6520
rect 44600 6508 44606 6520
rect 172514 6508 172520 6520
rect 44600 6480 172520 6508
rect 44600 6468 44606 6480
rect 172514 6468 172520 6480
rect 172572 6468 172578 6520
rect 344830 6468 344836 6520
rect 344888 6508 344894 6520
rect 469122 6508 469128 6520
rect 344888 6480 469128 6508
rect 344888 6468 344894 6480
rect 469122 6468 469128 6480
rect 469180 6468 469186 6520
rect 40954 6400 40960 6452
rect 41012 6440 41018 6452
rect 171226 6440 171232 6452
rect 41012 6412 171232 6440
rect 41012 6400 41018 6412
rect 171226 6400 171232 6412
rect 171284 6400 171290 6452
rect 178954 6400 178960 6452
rect 179012 6440 179018 6452
rect 226426 6440 226432 6452
rect 179012 6412 226432 6440
rect 179012 6400 179018 6412
rect 226426 6400 226432 6412
rect 226484 6400 226490 6452
rect 346302 6400 346308 6452
rect 346360 6440 346366 6452
rect 472710 6440 472716 6452
rect 346360 6412 472716 6440
rect 346360 6400 346366 6412
rect 472710 6400 472716 6412
rect 472768 6400 472774 6452
rect 37366 6332 37372 6384
rect 37424 6372 37430 6384
rect 169846 6372 169852 6384
rect 37424 6344 169852 6372
rect 37424 6332 37430 6344
rect 169846 6332 169852 6344
rect 169904 6332 169910 6384
rect 175366 6332 175372 6384
rect 175424 6372 175430 6384
rect 225046 6372 225052 6384
rect 175424 6344 225052 6372
rect 175424 6332 175430 6344
rect 225046 6332 225052 6344
rect 225104 6332 225110 6384
rect 347590 6332 347596 6384
rect 347648 6372 347654 6384
rect 476298 6372 476304 6384
rect 347648 6344 476304 6372
rect 347648 6332 347654 6344
rect 476298 6332 476304 6344
rect 476356 6332 476362 6384
rect 33870 6264 33876 6316
rect 33928 6304 33934 6316
rect 168466 6304 168472 6316
rect 33928 6276 168472 6304
rect 33928 6264 33934 6276
rect 168466 6264 168472 6276
rect 168524 6264 168530 6316
rect 171778 6264 171784 6316
rect 171836 6304 171842 6316
rect 223666 6304 223672 6316
rect 171836 6276 223672 6304
rect 171836 6264 171842 6276
rect 223666 6264 223672 6276
rect 223724 6264 223730 6316
rect 349062 6264 349068 6316
rect 349120 6304 349126 6316
rect 479886 6304 479892 6316
rect 349120 6276 479892 6304
rect 349120 6264 349126 6276
rect 479886 6264 479892 6276
rect 479944 6264 479950 6316
rect 8846 6196 8852 6248
rect 8904 6236 8910 6248
rect 157426 6236 157432 6248
rect 8904 6208 157432 6236
rect 8904 6196 8910 6208
rect 157426 6196 157432 6208
rect 157484 6196 157490 6248
rect 161106 6196 161112 6248
rect 161164 6236 161170 6248
rect 219434 6236 219440 6248
rect 161164 6208 219440 6236
rect 161164 6196 161170 6208
rect 219434 6196 219440 6208
rect 219492 6196 219498 6248
rect 277210 6196 277216 6248
rect 277268 6236 277274 6248
rect 302602 6236 302608 6248
rect 277268 6208 302608 6236
rect 277268 6196 277274 6208
rect 302602 6196 302608 6208
rect 302660 6196 302666 6248
rect 350350 6196 350356 6248
rect 350408 6236 350414 6248
rect 484578 6236 484584 6248
rect 350408 6208 484584 6236
rect 350408 6196 350414 6208
rect 484578 6196 484584 6208
rect 484636 6196 484642 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 156138 6168 156144 6180
rect 4120 6140 156144 6168
rect 4120 6128 4126 6140
rect 156138 6128 156144 6140
rect 156196 6128 156202 6180
rect 157518 6128 157524 6180
rect 157576 6168 157582 6180
rect 218146 6168 218152 6180
rect 157576 6140 218152 6168
rect 157576 6128 157582 6140
rect 218146 6128 218152 6140
rect 218204 6128 218210 6180
rect 272978 6128 272984 6180
rect 273036 6168 273042 6180
rect 273036 6140 287100 6168
rect 273036 6128 273042 6140
rect 136082 6060 136088 6112
rect 136140 6100 136146 6112
rect 210050 6100 210056 6112
rect 136140 6072 210056 6100
rect 136140 6060 136146 6072
rect 210050 6060 210056 6072
rect 210108 6060 210114 6112
rect 139670 5992 139676 6044
rect 139728 6032 139734 6044
rect 211338 6032 211344 6044
rect 139728 6004 211344 6032
rect 139728 5992 139734 6004
rect 211338 5992 211344 6004
rect 211396 5992 211402 6044
rect 287072 6032 287100 6140
rect 290458 6128 290464 6180
rect 290516 6168 290522 6180
rect 319254 6168 319260 6180
rect 290516 6140 319260 6168
rect 290516 6128 290522 6140
rect 319254 6128 319260 6140
rect 319312 6128 319318 6180
rect 351822 6128 351828 6180
rect 351880 6168 351886 6180
rect 488166 6168 488172 6180
rect 351880 6140 488172 6168
rect 351880 6128 351886 6140
rect 488166 6128 488172 6140
rect 488224 6128 488230 6180
rect 335262 6060 335268 6112
rect 335320 6100 335326 6112
rect 447778 6100 447784 6112
rect 335320 6072 447784 6100
rect 335320 6060 335326 6072
rect 447778 6060 447784 6072
rect 447836 6060 447842 6112
rect 290734 6032 290740 6044
rect 287072 6004 290740 6032
rect 290734 5992 290740 6004
rect 290792 5992 290798 6044
rect 333790 5992 333796 6044
rect 333848 6032 333854 6044
rect 444190 6032 444196 6044
rect 333848 6004 444196 6032
rect 333848 5992 333854 6004
rect 444190 5992 444196 6004
rect 444248 5992 444254 6044
rect 143258 5924 143264 5976
rect 143316 5964 143322 5976
rect 212534 5964 212540 5976
rect 143316 5936 212540 5964
rect 143316 5924 143322 5936
rect 212534 5924 212540 5936
rect 212592 5924 212598 5976
rect 332502 5924 332508 5976
rect 332560 5964 332566 5976
rect 440602 5964 440608 5976
rect 332560 5936 440608 5964
rect 332560 5924 332566 5936
rect 440602 5924 440608 5936
rect 440660 5924 440666 5976
rect 146846 5856 146852 5908
rect 146904 5896 146910 5908
rect 213914 5896 213920 5908
rect 146904 5868 213920 5896
rect 146904 5856 146910 5868
rect 213914 5856 213920 5868
rect 213972 5856 213978 5908
rect 331030 5856 331036 5908
rect 331088 5896 331094 5908
rect 437014 5896 437020 5908
rect 331088 5868 437020 5896
rect 331088 5856 331094 5868
rect 437014 5856 437020 5868
rect 437072 5856 437078 5908
rect 150434 5788 150440 5840
rect 150492 5828 150498 5840
rect 215478 5828 215484 5840
rect 150492 5800 215484 5828
rect 150492 5788 150498 5800
rect 215478 5788 215484 5800
rect 215536 5788 215542 5840
rect 222197 5831 222255 5837
rect 222197 5797 222209 5831
rect 222243 5828 222255 5831
rect 230474 5828 230480 5840
rect 222243 5800 230480 5828
rect 222243 5797 222255 5800
rect 222197 5791 222255 5797
rect 230474 5788 230480 5800
rect 230532 5788 230538 5840
rect 329742 5788 329748 5840
rect 329800 5828 329806 5840
rect 433518 5828 433524 5840
rect 329800 5800 433524 5828
rect 329800 5788 329806 5800
rect 433518 5788 433524 5800
rect 433576 5788 433582 5840
rect 153930 5720 153936 5772
rect 153988 5760 153994 5772
rect 216766 5760 216772 5772
rect 153988 5732 216772 5760
rect 153988 5720 153994 5732
rect 216766 5720 216772 5732
rect 216824 5720 216830 5772
rect 328270 5720 328276 5772
rect 328328 5760 328334 5772
rect 429930 5760 429936 5772
rect 328328 5732 429936 5760
rect 328328 5720 328334 5732
rect 429930 5720 429936 5732
rect 429988 5720 429994 5772
rect 164694 5652 164700 5704
rect 164752 5692 164758 5704
rect 220906 5692 220912 5704
rect 164752 5664 220912 5692
rect 164752 5652 164758 5664
rect 220906 5652 220912 5664
rect 220964 5652 220970 5704
rect 326982 5652 326988 5704
rect 327040 5692 327046 5704
rect 426342 5692 426348 5704
rect 327040 5664 426348 5692
rect 327040 5652 327046 5664
rect 426342 5652 426348 5664
rect 426400 5652 426406 5704
rect 168190 5584 168196 5636
rect 168248 5624 168254 5636
rect 222286 5624 222292 5636
rect 168248 5596 222292 5624
rect 168248 5584 168254 5596
rect 222286 5584 222292 5596
rect 222344 5584 222350 5636
rect 325510 5584 325516 5636
rect 325568 5624 325574 5636
rect 422754 5624 422760 5636
rect 325568 5596 422760 5624
rect 325568 5584 325574 5596
rect 422754 5584 422760 5596
rect 422812 5584 422818 5636
rect 287698 5516 287704 5568
rect 287756 5556 287762 5568
rect 294322 5556 294328 5568
rect 287756 5528 294328 5556
rect 287756 5516 287762 5528
rect 294322 5516 294328 5528
rect 294380 5516 294386 5568
rect 51626 5448 51632 5500
rect 51684 5488 51690 5500
rect 175274 5488 175280 5500
rect 51684 5460 175280 5488
rect 51684 5448 51690 5460
rect 175274 5448 175280 5460
rect 175332 5448 175338 5500
rect 197998 5448 198004 5500
rect 198056 5488 198062 5500
rect 234706 5488 234712 5500
rect 198056 5460 234712 5488
rect 198056 5448 198062 5460
rect 234706 5448 234712 5460
rect 234764 5448 234770 5500
rect 296438 5448 296444 5500
rect 296496 5488 296502 5500
rect 351362 5488 351368 5500
rect 296496 5460 351368 5488
rect 296496 5448 296502 5460
rect 351362 5448 351368 5460
rect 351420 5448 351426 5500
rect 375190 5448 375196 5500
rect 375248 5488 375254 5500
rect 544102 5488 544108 5500
rect 375248 5460 544108 5488
rect 375248 5448 375254 5460
rect 544102 5448 544108 5460
rect 544160 5448 544166 5500
rect 48130 5380 48136 5432
rect 48188 5420 48194 5432
rect 173986 5420 173992 5432
rect 48188 5392 173992 5420
rect 48188 5380 48194 5392
rect 173986 5380 173992 5392
rect 174044 5380 174050 5432
rect 190822 5380 190828 5432
rect 190880 5420 190886 5432
rect 230566 5420 230572 5432
rect 190880 5392 230572 5420
rect 190880 5380 190886 5392
rect 230566 5380 230572 5392
rect 230624 5380 230630 5432
rect 297818 5380 297824 5432
rect 297876 5420 297882 5432
rect 354950 5420 354956 5432
rect 297876 5392 354956 5420
rect 297876 5380 297882 5392
rect 354950 5380 354956 5392
rect 355008 5380 355014 5432
rect 376570 5380 376576 5432
rect 376628 5420 376634 5432
rect 547690 5420 547696 5432
rect 376628 5392 547696 5420
rect 376628 5380 376634 5392
rect 547690 5380 547696 5392
rect 547748 5380 547754 5432
rect 30282 5312 30288 5364
rect 30340 5352 30346 5364
rect 167178 5352 167184 5364
rect 30340 5324 167184 5352
rect 30340 5312 30346 5324
rect 167178 5312 167184 5324
rect 167236 5312 167242 5364
rect 194502 5312 194508 5364
rect 194560 5352 194566 5364
rect 233326 5352 233332 5364
rect 194560 5324 233332 5352
rect 194560 5312 194566 5324
rect 233326 5312 233332 5324
rect 233384 5312 233390 5364
rect 299290 5312 299296 5364
rect 299348 5352 299354 5364
rect 358538 5352 358544 5364
rect 299348 5324 358544 5352
rect 299348 5312 299354 5324
rect 358538 5312 358544 5324
rect 358596 5312 358602 5364
rect 377950 5312 377956 5364
rect 378008 5352 378014 5364
rect 551186 5352 551192 5364
rect 378008 5324 551192 5352
rect 378008 5312 378014 5324
rect 551186 5312 551192 5324
rect 551244 5312 551250 5364
rect 26694 5244 26700 5296
rect 26752 5284 26758 5296
rect 165706 5284 165712 5296
rect 26752 5256 165712 5284
rect 26752 5244 26758 5256
rect 165706 5244 165712 5256
rect 165764 5244 165770 5296
rect 181346 5244 181352 5296
rect 181404 5284 181410 5296
rect 227714 5284 227720 5296
rect 181404 5256 227720 5284
rect 181404 5244 181410 5256
rect 227714 5244 227720 5256
rect 227772 5244 227778 5296
rect 300670 5244 300676 5296
rect 300728 5284 300734 5296
rect 362126 5284 362132 5296
rect 300728 5256 362132 5284
rect 300728 5244 300734 5256
rect 362126 5244 362132 5256
rect 362184 5244 362190 5296
rect 379330 5244 379336 5296
rect 379388 5284 379394 5296
rect 554774 5284 554780 5296
rect 379388 5256 554780 5284
rect 379388 5244 379394 5256
rect 554774 5244 554780 5256
rect 554832 5244 554838 5296
rect 21910 5176 21916 5228
rect 21968 5216 21974 5228
rect 163130 5216 163136 5228
rect 21968 5188 163136 5216
rect 21968 5176 21974 5188
rect 163130 5176 163136 5188
rect 163188 5176 163194 5228
rect 177758 5176 177764 5228
rect 177816 5216 177822 5228
rect 226334 5216 226340 5228
rect 177816 5188 226340 5216
rect 177816 5176 177822 5188
rect 226334 5176 226340 5188
rect 226392 5176 226398 5228
rect 303430 5176 303436 5228
rect 303488 5216 303494 5228
rect 365714 5216 365720 5228
rect 303488 5188 365720 5216
rect 303488 5176 303494 5188
rect 365714 5176 365720 5188
rect 365772 5176 365778 5228
rect 380710 5176 380716 5228
rect 380768 5216 380774 5228
rect 558362 5216 558368 5228
rect 380768 5188 558368 5216
rect 380768 5176 380774 5188
rect 558362 5176 558368 5188
rect 558420 5176 558426 5228
rect 17218 5108 17224 5160
rect 17276 5148 17282 5160
rect 161474 5148 161480 5160
rect 17276 5120 161480 5148
rect 17276 5108 17282 5120
rect 161474 5108 161480 5120
rect 161532 5108 161538 5160
rect 174170 5108 174176 5160
rect 174228 5148 174234 5160
rect 224954 5148 224960 5160
rect 174228 5120 224960 5148
rect 174228 5108 174234 5120
rect 224954 5108 224960 5120
rect 225012 5108 225018 5160
rect 304810 5108 304816 5160
rect 304868 5148 304874 5160
rect 369210 5148 369216 5160
rect 304868 5120 369216 5148
rect 304868 5108 304874 5120
rect 369210 5108 369216 5120
rect 369268 5108 369274 5160
rect 382090 5108 382096 5160
rect 382148 5148 382154 5160
rect 561950 5148 561956 5160
rect 382148 5120 561956 5148
rect 382148 5108 382154 5120
rect 561950 5108 561956 5120
rect 562008 5108 562014 5160
rect 12434 5040 12440 5092
rect 12492 5080 12498 5092
rect 158806 5080 158812 5092
rect 12492 5052 158812 5080
rect 12492 5040 12498 5052
rect 158806 5040 158812 5052
rect 158864 5040 158870 5092
rect 170582 5040 170588 5092
rect 170640 5080 170646 5092
rect 223574 5080 223580 5092
rect 170640 5052 223580 5080
rect 170640 5040 170646 5052
rect 223574 5040 223580 5052
rect 223632 5040 223638 5092
rect 306190 5040 306196 5092
rect 306248 5080 306254 5092
rect 372798 5080 372804 5092
rect 306248 5052 372804 5080
rect 306248 5040 306254 5052
rect 372798 5040 372804 5052
rect 372856 5040 372862 5092
rect 383562 5040 383568 5092
rect 383620 5080 383626 5092
rect 565538 5080 565544 5092
rect 383620 5052 565544 5080
rect 383620 5040 383626 5052
rect 565538 5040 565544 5052
rect 565596 5040 565602 5092
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 157702 5012 157708 5024
rect 7708 4984 157708 5012
rect 7708 4972 7714 4984
rect 157702 4972 157708 4984
rect 157760 4972 157766 5024
rect 167086 4972 167092 5024
rect 167144 5012 167150 5024
rect 222194 5012 222200 5024
rect 167144 4984 222200 5012
rect 167144 4972 167150 4984
rect 222194 4972 222200 4984
rect 222252 4972 222258 5024
rect 307662 4972 307668 5024
rect 307720 5012 307726 5024
rect 376386 5012 376392 5024
rect 307720 4984 376392 5012
rect 307720 4972 307726 4984
rect 376386 4972 376392 4984
rect 376444 4972 376450 5024
rect 384850 4972 384856 5024
rect 384908 5012 384914 5024
rect 569034 5012 569040 5024
rect 384908 4984 569040 5012
rect 384908 4972 384914 4984
rect 569034 4972 569040 4984
rect 569092 4972 569098 5024
rect 1670 4904 1676 4956
rect 1728 4944 1734 4956
rect 154574 4944 154580 4956
rect 1728 4916 154580 4944
rect 1728 4904 1734 4916
rect 154574 4904 154580 4916
rect 154632 4904 154638 4956
rect 163498 4904 163504 4956
rect 163556 4944 163562 4956
rect 220814 4944 220820 4956
rect 163556 4916 220820 4944
rect 163556 4904 163562 4916
rect 220814 4904 220820 4916
rect 220872 4904 220878 4956
rect 308950 4904 308956 4956
rect 309008 4944 309014 4956
rect 379974 4944 379980 4956
rect 309008 4916 379980 4944
rect 309008 4904 309014 4916
rect 379974 4904 379980 4916
rect 380032 4904 380038 4956
rect 386230 4904 386236 4956
rect 386288 4944 386294 4956
rect 572622 4944 572628 4956
rect 386288 4916 572628 4944
rect 386288 4904 386294 4916
rect 572622 4904 572628 4916
rect 572680 4904 572686 4956
rect 2866 4836 2872 4888
rect 2924 4876 2930 4888
rect 156046 4876 156052 4888
rect 2924 4848 156052 4876
rect 2924 4836 2930 4848
rect 156046 4836 156052 4848
rect 156104 4836 156110 4888
rect 158714 4836 158720 4888
rect 158772 4876 158778 4888
rect 218054 4876 218060 4888
rect 158772 4848 218060 4876
rect 158772 4836 158778 4848
rect 218054 4836 218060 4848
rect 218112 4836 218118 4888
rect 310422 4836 310428 4888
rect 310480 4876 310486 4888
rect 383562 4876 383568 4888
rect 310480 4848 383568 4876
rect 310480 4836 310486 4848
rect 383562 4836 383568 4848
rect 383620 4836 383626 4888
rect 387610 4836 387616 4888
rect 387668 4876 387674 4888
rect 576210 4876 576216 4888
rect 387668 4848 576216 4876
rect 387668 4836 387674 4848
rect 576210 4836 576216 4848
rect 576268 4836 576274 4888
rect 566 4768 572 4820
rect 624 4808 630 4820
rect 154666 4808 154672 4820
rect 624 4780 154672 4808
rect 624 4768 630 4780
rect 154666 4768 154672 4780
rect 154724 4768 154730 4820
rect 155126 4768 155132 4820
rect 155184 4808 155190 4820
rect 216950 4808 216956 4820
rect 155184 4780 216956 4808
rect 155184 4768 155190 4780
rect 216950 4768 216956 4780
rect 217008 4768 217014 4820
rect 230477 4811 230535 4817
rect 230477 4777 230489 4811
rect 230523 4808 230535 4811
rect 233418 4808 233424 4820
rect 230523 4780 233424 4808
rect 230523 4777 230535 4780
rect 230477 4771 230535 4777
rect 233418 4768 233424 4780
rect 233476 4768 233482 4820
rect 270218 4768 270224 4820
rect 270276 4808 270282 4820
rect 283650 4808 283656 4820
rect 270276 4780 283656 4808
rect 270276 4768 270282 4780
rect 283650 4768 283656 4780
rect 283708 4768 283714 4820
rect 311710 4768 311716 4820
rect 311768 4808 311774 4820
rect 387058 4808 387064 4820
rect 311768 4780 387064 4808
rect 311768 4768 311774 4780
rect 387058 4768 387064 4780
rect 387116 4768 387122 4820
rect 388990 4768 388996 4820
rect 389048 4808 389054 4820
rect 579798 4808 579804 4820
rect 389048 4780 579804 4808
rect 389048 4768 389054 4780
rect 579798 4768 579804 4780
rect 579856 4768 579862 4820
rect 55214 4700 55220 4752
rect 55272 4740 55278 4752
rect 176654 4740 176660 4752
rect 55272 4712 176660 4740
rect 55272 4700 55278 4712
rect 176654 4700 176660 4712
rect 176712 4700 176718 4752
rect 297910 4700 297916 4752
rect 297968 4740 297974 4752
rect 352558 4740 352564 4752
rect 297968 4712 352564 4740
rect 297968 4700 297974 4712
rect 352558 4700 352564 4712
rect 352616 4700 352622 4752
rect 371142 4700 371148 4752
rect 371200 4740 371206 4752
rect 536926 4740 536932 4752
rect 371200 4712 536932 4740
rect 371200 4700 371206 4712
rect 536926 4700 536932 4712
rect 536984 4700 536990 4752
rect 58802 4632 58808 4684
rect 58860 4672 58866 4684
rect 178034 4672 178040 4684
rect 58860 4644 178040 4672
rect 58860 4632 58866 4644
rect 178034 4632 178040 4644
rect 178092 4632 178098 4684
rect 295150 4632 295156 4684
rect 295208 4672 295214 4684
rect 347866 4672 347872 4684
rect 295208 4644 347872 4672
rect 295208 4632 295214 4644
rect 347866 4632 347872 4644
rect 347924 4632 347930 4684
rect 373902 4632 373908 4684
rect 373960 4672 373966 4684
rect 540514 4672 540520 4684
rect 373960 4644 540520 4672
rect 373960 4632 373966 4644
rect 540514 4632 540520 4644
rect 540572 4632 540578 4684
rect 62390 4564 62396 4616
rect 62448 4604 62454 4616
rect 179414 4604 179420 4616
rect 62448 4576 179420 4604
rect 62448 4564 62454 4576
rect 179414 4564 179420 4576
rect 179472 4564 179478 4616
rect 296530 4564 296536 4616
rect 296588 4604 296594 4616
rect 349062 4604 349068 4616
rect 296588 4576 349068 4604
rect 296588 4564 296594 4576
rect 349062 4564 349068 4576
rect 349120 4564 349126 4616
rect 369762 4564 369768 4616
rect 369820 4604 369826 4616
rect 533430 4604 533436 4616
rect 369820 4576 533436 4604
rect 369820 4564 369826 4576
rect 533430 4564 533436 4576
rect 533488 4564 533494 4616
rect 65978 4496 65984 4548
rect 66036 4536 66042 4548
rect 180886 4536 180892 4548
rect 66036 4508 180892 4536
rect 66036 4496 66042 4508
rect 180886 4496 180892 4508
rect 180944 4496 180950 4548
rect 293678 4496 293684 4548
rect 293736 4536 293742 4548
rect 344278 4536 344284 4548
rect 293736 4508 344284 4536
rect 293736 4496 293742 4508
rect 344278 4496 344284 4508
rect 344336 4496 344342 4548
rect 368382 4496 368388 4548
rect 368440 4536 368446 4548
rect 529842 4536 529848 4548
rect 368440 4508 529848 4536
rect 368440 4496 368446 4508
rect 529842 4496 529848 4508
rect 529900 4496 529906 4548
rect 69474 4428 69480 4480
rect 69532 4468 69538 4480
rect 182266 4468 182272 4480
rect 69532 4440 182272 4468
rect 69532 4428 69538 4440
rect 182266 4428 182272 4440
rect 182324 4428 182330 4480
rect 295058 4428 295064 4480
rect 295116 4468 295122 4480
rect 345474 4468 345480 4480
rect 295116 4440 345480 4468
rect 295116 4428 295122 4440
rect 345474 4428 345480 4440
rect 345532 4428 345538 4480
rect 367002 4428 367008 4480
rect 367060 4468 367066 4480
rect 526254 4468 526260 4480
rect 367060 4440 526260 4468
rect 367060 4428 367066 4440
rect 526254 4428 526260 4440
rect 526312 4428 526318 4480
rect 73062 4360 73068 4412
rect 73120 4400 73126 4412
rect 183646 4400 183652 4412
rect 73120 4372 183652 4400
rect 73120 4360 73126 4372
rect 183646 4360 183652 4372
rect 183704 4360 183710 4412
rect 293770 4360 293776 4412
rect 293828 4400 293834 4412
rect 341886 4400 341892 4412
rect 293828 4372 341892 4400
rect 293828 4360 293834 4372
rect 341886 4360 341892 4372
rect 341944 4360 341950 4412
rect 365622 4360 365628 4412
rect 365680 4400 365686 4412
rect 522666 4400 522672 4412
rect 365680 4372 522672 4400
rect 365680 4360 365686 4372
rect 522666 4360 522672 4372
rect 522724 4360 522730 4412
rect 76650 4292 76656 4344
rect 76708 4332 76714 4344
rect 185121 4335 185179 4341
rect 185121 4332 185133 4335
rect 76708 4304 185133 4332
rect 76708 4292 76714 4304
rect 185121 4301 185133 4304
rect 185167 4301 185179 4335
rect 185121 4295 185179 4301
rect 292390 4292 292396 4344
rect 292448 4332 292454 4344
rect 338298 4332 338304 4344
rect 292448 4304 338304 4332
rect 292448 4292 292454 4304
rect 338298 4292 338304 4304
rect 338356 4292 338362 4344
rect 364242 4292 364248 4344
rect 364300 4332 364306 4344
rect 519078 4332 519084 4344
rect 364300 4304 519084 4332
rect 364300 4292 364306 4304
rect 519078 4292 519084 4304
rect 519136 4292 519142 4344
rect 80238 4224 80244 4276
rect 80296 4264 80302 4276
rect 186406 4264 186412 4276
rect 80296 4236 186412 4264
rect 80296 4224 80302 4236
rect 186406 4224 186412 4236
rect 186464 4224 186470 4276
rect 289630 4224 289636 4276
rect 289688 4264 289694 4276
rect 334710 4264 334716 4276
rect 289688 4236 334716 4264
rect 289688 4224 289694 4236
rect 334710 4224 334716 4236
rect 334768 4224 334774 4276
rect 362862 4224 362868 4276
rect 362920 4264 362926 4276
rect 515582 4264 515588 4276
rect 362920 4236 515588 4264
rect 362920 4224 362926 4236
rect 515582 4224 515588 4236
rect 515640 4224 515646 4276
rect 140866 4156 140872 4208
rect 140924 4196 140930 4208
rect 142062 4196 142068 4208
rect 140924 4168 142068 4196
rect 140924 4156 140930 4168
rect 142062 4156 142068 4168
rect 142120 4156 142126 4208
rect 222856 4168 223620 4196
rect 14826 4088 14832 4140
rect 14884 4128 14890 4140
rect 18598 4128 18604 4140
rect 14884 4100 18604 4128
rect 14884 4088 14890 4100
rect 18598 4088 18604 4100
rect 18656 4088 18662 4140
rect 93765 4131 93823 4137
rect 93765 4097 93777 4131
rect 93811 4128 93823 4131
rect 187694 4128 187700 4140
rect 93811 4100 187700 4128
rect 93811 4097 93823 4100
rect 93765 4091 93823 4097
rect 187694 4088 187700 4100
rect 187752 4088 187758 4140
rect 188430 4088 188436 4140
rect 188488 4128 188494 4140
rect 188982 4128 188988 4140
rect 188488 4100 188988 4128
rect 188488 4088 188494 4100
rect 188982 4088 188988 4100
rect 189040 4088 189046 4140
rect 199194 4088 199200 4140
rect 199252 4128 199258 4140
rect 200022 4128 200028 4140
rect 199252 4100 200028 4128
rect 199252 4088 199258 4100
rect 200022 4088 200028 4100
rect 200080 4088 200086 4140
rect 200390 4088 200396 4140
rect 200448 4128 200454 4140
rect 201402 4128 201408 4140
rect 200448 4100 201408 4128
rect 200448 4088 200454 4100
rect 201402 4088 201408 4100
rect 201460 4088 201466 4140
rect 206278 4088 206284 4140
rect 206336 4128 206342 4140
rect 206922 4128 206928 4140
rect 206336 4100 206928 4128
rect 206336 4088 206342 4100
rect 206922 4088 206928 4100
rect 206980 4088 206986 4140
rect 215846 4088 215852 4140
rect 215904 4128 215910 4140
rect 216582 4128 216588 4140
rect 215904 4100 216588 4128
rect 215904 4088 215910 4100
rect 216582 4088 216588 4100
rect 216640 4088 216646 4140
rect 217042 4088 217048 4140
rect 217100 4128 217106 4140
rect 217962 4128 217968 4140
rect 217100 4100 217968 4128
rect 217100 4088 217106 4100
rect 217962 4088 217968 4100
rect 218020 4088 218026 4140
rect 218146 4088 218152 4140
rect 218204 4128 218210 4140
rect 222856 4128 222884 4168
rect 218204 4100 222884 4128
rect 218204 4088 218210 4100
rect 222930 4088 222936 4140
rect 222988 4128 222994 4140
rect 223482 4128 223488 4140
rect 222988 4100 223488 4128
rect 222988 4088 222994 4100
rect 223482 4088 223488 4100
rect 223540 4088 223546 4140
rect 223592 4128 223620 4168
rect 234709 4131 234767 4137
rect 234709 4128 234721 4131
rect 223592 4100 234721 4128
rect 234709 4097 234721 4100
rect 234755 4097 234767 4131
rect 234709 4091 234767 4097
rect 234798 4088 234804 4140
rect 234856 4128 234862 4140
rect 235902 4128 235908 4140
rect 234856 4100 235908 4128
rect 234856 4088 234862 4100
rect 235902 4088 235908 4100
rect 235960 4088 235966 4140
rect 240778 4088 240784 4140
rect 240836 4128 240842 4140
rect 241422 4128 241428 4140
rect 240836 4100 241428 4128
rect 240836 4088 240842 4100
rect 241422 4088 241428 4100
rect 241480 4088 241486 4140
rect 244274 4128 244280 4140
rect 241532 4100 244280 4128
rect 82630 4020 82636 4072
rect 82688 4060 82694 4072
rect 84749 4063 84807 4069
rect 84749 4060 84761 4063
rect 82688 4032 84761 4060
rect 82688 4020 82694 4032
rect 84749 4029 84761 4032
rect 84795 4029 84807 4063
rect 84749 4023 84807 4029
rect 84841 4063 84899 4069
rect 84841 4029 84853 4063
rect 84887 4060 84899 4063
rect 186314 4060 186320 4072
rect 84887 4032 186320 4060
rect 84887 4029 84899 4032
rect 84841 4023 84899 4029
rect 186314 4020 186320 4032
rect 186372 4020 186378 4072
rect 221734 4020 221740 4072
rect 221792 4060 221798 4072
rect 241532 4060 241560 4100
rect 244274 4088 244280 4100
rect 244332 4088 244338 4140
rect 244366 4088 244372 4140
rect 244424 4128 244430 4140
rect 245562 4128 245568 4140
rect 244424 4100 245568 4128
rect 244424 4088 244430 4100
rect 245562 4088 245568 4100
rect 245620 4088 245626 4140
rect 257430 4088 257436 4140
rect 257488 4128 257494 4140
rect 257982 4128 257988 4140
rect 257488 4100 257988 4128
rect 257488 4088 257494 4100
rect 257982 4088 257988 4100
rect 258040 4088 258046 4140
rect 258166 4088 258172 4140
rect 258224 4128 258230 4140
rect 258626 4128 258632 4140
rect 258224 4100 258632 4128
rect 258224 4088 258230 4100
rect 258626 4088 258632 4100
rect 258684 4088 258690 4140
rect 262122 4088 262128 4140
rect 262180 4128 262186 4140
rect 263410 4128 263416 4140
rect 262180 4100 263416 4128
rect 262180 4088 262186 4100
rect 263410 4088 263416 4100
rect 263468 4088 263474 4140
rect 270310 4088 270316 4140
rect 270368 4128 270374 4140
rect 284754 4128 284760 4140
rect 270368 4100 284760 4128
rect 270368 4088 270374 4100
rect 284754 4088 284760 4100
rect 284812 4088 284818 4140
rect 289722 4088 289728 4140
rect 289780 4128 289786 4140
rect 332410 4128 332416 4140
rect 289780 4100 332416 4128
rect 289780 4088 289786 4100
rect 332410 4088 332416 4100
rect 332468 4088 332474 4140
rect 339402 4088 339408 4140
rect 339460 4128 339466 4140
rect 457254 4128 457260 4140
rect 339460 4100 457260 4128
rect 339460 4088 339466 4100
rect 457254 4088 457260 4100
rect 457312 4088 457318 4140
rect 221792 4032 241560 4060
rect 221792 4020 221798 4032
rect 243170 4020 243176 4072
rect 243228 4060 243234 4072
rect 244918 4060 244924 4072
rect 243228 4032 244924 4060
rect 243228 4020 243234 4032
rect 244918 4020 244924 4032
rect 244976 4020 244982 4072
rect 260742 4020 260748 4072
rect 260800 4060 260806 4072
rect 262214 4060 262220 4072
rect 260800 4032 262220 4060
rect 260800 4020 260806 4032
rect 262214 4020 262220 4032
rect 262272 4020 262278 4072
rect 270402 4020 270408 4072
rect 270460 4060 270466 4072
rect 285950 4060 285956 4072
rect 270460 4032 285956 4060
rect 270460 4020 270466 4032
rect 285950 4020 285956 4032
rect 286008 4020 286014 4072
rect 291102 4020 291108 4072
rect 291160 4060 291166 4072
rect 335906 4060 335912 4072
rect 291160 4032 335912 4060
rect 291160 4020 291166 4032
rect 335906 4020 335912 4032
rect 335964 4020 335970 4072
rect 342162 4020 342168 4072
rect 342220 4060 342226 4072
rect 464430 4060 464436 4072
rect 342220 4032 464436 4060
rect 342220 4020 342226 4032
rect 464430 4020 464436 4032
rect 464488 4020 464494 4072
rect 75454 3952 75460 4004
rect 75512 3992 75518 4004
rect 75512 3964 180012 3992
rect 75512 3952 75518 3964
rect 71866 3884 71872 3936
rect 71924 3924 71930 3936
rect 71924 3896 176700 3924
rect 71924 3884 71930 3896
rect 68278 3816 68284 3868
rect 68336 3856 68342 3868
rect 170585 3859 170643 3865
rect 170585 3856 170597 3859
rect 68336 3828 170597 3856
rect 68336 3816 68342 3828
rect 170585 3825 170597 3828
rect 170631 3825 170643 3859
rect 170585 3819 170643 3825
rect 172974 3816 172980 3868
rect 173032 3856 173038 3868
rect 173802 3856 173808 3868
rect 173032 3828 173808 3856
rect 173032 3816 173038 3828
rect 173802 3816 173808 3828
rect 173860 3816 173866 3868
rect 64782 3748 64788 3800
rect 64840 3788 64846 3800
rect 166997 3791 167055 3797
rect 166997 3788 167009 3791
rect 64840 3760 167009 3788
rect 64840 3748 64846 3760
rect 166997 3757 167009 3760
rect 167043 3757 167055 3791
rect 176672 3788 176700 3896
rect 179984 3856 180012 3964
rect 180150 3952 180156 4004
rect 180208 3992 180214 4004
rect 180702 3992 180708 4004
rect 180208 3964 180708 3992
rect 180208 3952 180214 3964
rect 180702 3952 180708 3964
rect 180760 3952 180766 4004
rect 182542 3952 182548 4004
rect 182600 3992 182606 4004
rect 183462 3992 183468 4004
rect 182600 3964 183468 3992
rect 182600 3952 182606 3964
rect 183462 3952 183468 3964
rect 183520 3952 183526 4004
rect 208670 3952 208676 4004
rect 208728 3992 208734 4004
rect 220081 3995 220139 4001
rect 220081 3992 220093 3995
rect 208728 3964 220093 3992
rect 208728 3952 208734 3964
rect 220081 3961 220093 3964
rect 220127 3961 220139 3995
rect 220081 3955 220139 3961
rect 220538 3952 220544 4004
rect 220596 3992 220602 4004
rect 234617 3995 234675 4001
rect 234617 3992 234629 3995
rect 220596 3964 234629 3992
rect 220596 3952 220602 3964
rect 234617 3961 234629 3964
rect 234663 3961 234675 3995
rect 234617 3955 234675 3961
rect 234709 3995 234767 4001
rect 234709 3961 234721 3995
rect 234755 3992 234767 3995
rect 241606 3992 241612 4004
rect 234755 3964 241612 3992
rect 234755 3961 234767 3964
rect 234709 3955 234767 3961
rect 241606 3952 241612 3964
rect 241664 3952 241670 4004
rect 266998 3952 267004 4004
rect 267056 3992 267062 4004
rect 270494 3992 270500 4004
rect 267056 3964 270500 3992
rect 267056 3952 267062 3964
rect 270494 3952 270500 3964
rect 270552 3952 270558 4004
rect 271690 3952 271696 4004
rect 271748 3992 271754 4004
rect 288342 3992 288348 4004
rect 271748 3964 288348 3992
rect 271748 3952 271754 3964
rect 288342 3952 288348 3964
rect 288400 3952 288406 4004
rect 292482 3952 292488 4004
rect 292540 3992 292546 4004
rect 339494 3992 339500 4004
rect 292540 3964 339500 3992
rect 292540 3952 292546 3964
rect 339494 3952 339500 3964
rect 339552 3952 339558 4004
rect 344922 3952 344928 4004
rect 344980 3992 344986 4004
rect 471514 3992 471520 4004
rect 344980 3964 471520 3992
rect 344980 3952 344986 3964
rect 471514 3952 471520 3964
rect 471572 3952 471578 4004
rect 214650 3884 214656 3936
rect 214708 3924 214714 3936
rect 226429 3927 226487 3933
rect 226429 3924 226441 3927
rect 214708 3896 226441 3924
rect 214708 3884 214714 3896
rect 226429 3893 226441 3896
rect 226475 3893 226487 3927
rect 226429 3887 226487 3893
rect 226518 3884 226524 3936
rect 226576 3924 226582 3936
rect 227622 3924 227628 3936
rect 226576 3896 227628 3924
rect 226576 3884 226582 3896
rect 227622 3884 227628 3896
rect 227680 3884 227686 3936
rect 240226 3924 240232 3936
rect 229664 3896 240232 3924
rect 184934 3856 184940 3868
rect 179984 3828 184940 3856
rect 184934 3816 184940 3828
rect 184992 3816 184998 3868
rect 209866 3816 209872 3868
rect 209924 3856 209930 3868
rect 229465 3859 229523 3865
rect 229465 3856 229477 3859
rect 209924 3828 229477 3856
rect 209924 3816 209930 3828
rect 229465 3825 229477 3828
rect 229511 3825 229523 3859
rect 229465 3819 229523 3825
rect 183554 3788 183560 3800
rect 176672 3760 183560 3788
rect 166997 3751 167055 3757
rect 183554 3748 183560 3760
rect 183612 3748 183618 3800
rect 211157 3791 211215 3797
rect 211157 3757 211169 3791
rect 211203 3788 211215 3791
rect 220725 3791 220783 3797
rect 220725 3788 220737 3791
rect 211203 3760 220737 3788
rect 211203 3757 211215 3760
rect 211157 3751 211215 3757
rect 220725 3757 220737 3760
rect 220771 3757 220783 3791
rect 220725 3751 220783 3757
rect 224865 3791 224923 3797
rect 224865 3757 224877 3791
rect 224911 3788 224923 3791
rect 229664 3788 229692 3896
rect 240226 3884 240232 3896
rect 240284 3884 240290 3936
rect 264238 3884 264244 3936
rect 264296 3924 264302 3936
rect 268102 3924 268108 3936
rect 264296 3896 268108 3924
rect 264296 3884 264302 3896
rect 268102 3884 268108 3896
rect 268160 3884 268166 3936
rect 271782 3884 271788 3936
rect 271840 3924 271846 3936
rect 289538 3924 289544 3936
rect 271840 3896 289544 3924
rect 271840 3884 271846 3896
rect 289538 3884 289544 3896
rect 289596 3884 289602 3936
rect 293862 3884 293868 3936
rect 293920 3924 293926 3936
rect 343082 3924 343088 3936
rect 293920 3896 343088 3924
rect 293920 3884 293926 3896
rect 343082 3884 343088 3896
rect 343140 3884 343146 3936
rect 347682 3884 347688 3936
rect 347740 3924 347746 3936
rect 478690 3924 478696 3936
rect 347740 3896 478696 3924
rect 347740 3884 347746 3896
rect 478690 3884 478696 3896
rect 478748 3884 478754 3936
rect 485774 3884 485780 3936
rect 485832 3924 485838 3936
rect 486970 3924 486976 3936
rect 485832 3896 486976 3924
rect 485832 3884 485838 3896
rect 486970 3884 486976 3896
rect 487028 3884 487034 3936
rect 494146 3884 494152 3936
rect 494204 3924 494210 3936
rect 495342 3924 495348 3936
rect 494204 3896 495348 3924
rect 494204 3884 494210 3896
rect 495342 3884 495348 3896
rect 495400 3884 495406 3936
rect 502426 3884 502432 3936
rect 502484 3924 502490 3936
rect 503622 3924 503628 3936
rect 502484 3896 503628 3924
rect 502484 3884 502490 3896
rect 503622 3884 503628 3896
rect 503680 3884 503686 3936
rect 229741 3859 229799 3865
rect 229741 3825 229753 3859
rect 229787 3856 229799 3859
rect 239030 3856 239036 3868
rect 229787 3828 239036 3856
rect 229787 3825 229799 3828
rect 229741 3819 229799 3825
rect 239030 3816 239036 3828
rect 239088 3816 239094 3868
rect 268838 3816 268844 3868
rect 268896 3856 268902 3868
rect 268896 3828 273024 3856
rect 268896 3816 268902 3828
rect 238846 3788 238852 3800
rect 224911 3760 229692 3788
rect 229756 3760 238852 3788
rect 224911 3757 224923 3760
rect 224865 3751 224923 3757
rect 46934 3680 46940 3732
rect 46992 3720 46998 3732
rect 173894 3720 173900 3732
rect 46992 3692 173900 3720
rect 46992 3680 46998 3692
rect 173894 3680 173900 3692
rect 173952 3680 173958 3732
rect 173989 3723 174047 3729
rect 173989 3689 174001 3723
rect 174035 3720 174047 3723
rect 180794 3720 180800 3732
rect 174035 3692 180800 3720
rect 174035 3689 174047 3692
rect 173989 3683 174047 3689
rect 180794 3680 180800 3692
rect 180852 3680 180858 3732
rect 220081 3723 220139 3729
rect 220081 3689 220093 3723
rect 220127 3720 220139 3723
rect 229756 3720 229784 3760
rect 238846 3748 238852 3760
rect 238904 3748 238910 3800
rect 264790 3748 264796 3800
rect 264848 3788 264854 3800
rect 271690 3788 271696 3800
rect 264848 3760 271696 3788
rect 264848 3748 264854 3760
rect 271690 3748 271696 3760
rect 271748 3748 271754 3800
rect 220127 3692 229784 3720
rect 220127 3689 220139 3692
rect 220081 3683 220139 3689
rect 230106 3680 230112 3732
rect 230164 3720 230170 3732
rect 231118 3720 231124 3732
rect 230164 3692 231124 3720
rect 230164 3680 230170 3692
rect 231118 3680 231124 3692
rect 231176 3680 231182 3732
rect 233694 3680 233700 3732
rect 233752 3720 233758 3732
rect 234522 3720 234528 3732
rect 233752 3692 234528 3720
rect 233752 3680 233758 3692
rect 234522 3680 234528 3692
rect 234580 3680 234586 3732
rect 234617 3723 234675 3729
rect 234617 3689 234629 3723
rect 234663 3720 234675 3723
rect 242894 3720 242900 3732
rect 234663 3692 242900 3720
rect 234663 3689 234675 3692
rect 234617 3683 234675 3689
rect 242894 3680 242900 3692
rect 242952 3680 242958 3732
rect 264882 3680 264888 3732
rect 264940 3720 264946 3732
rect 272886 3720 272892 3732
rect 264940 3692 272892 3720
rect 264940 3680 264946 3692
rect 272886 3680 272892 3692
rect 272944 3680 272950 3732
rect 272996 3720 273024 3828
rect 273070 3816 273076 3868
rect 273128 3856 273134 3868
rect 291930 3856 291936 3868
rect 273128 3828 291936 3856
rect 273128 3816 273134 3828
rect 291930 3816 291936 3828
rect 291988 3816 291994 3868
rect 295242 3816 295248 3868
rect 295300 3856 295306 3868
rect 346670 3856 346676 3868
rect 295300 3828 346676 3856
rect 295300 3816 295306 3828
rect 346670 3816 346676 3828
rect 346728 3816 346734 3868
rect 375282 3816 375288 3868
rect 375340 3856 375346 3868
rect 546494 3856 546500 3868
rect 375340 3828 546500 3856
rect 375340 3816 375346 3828
rect 546494 3816 546500 3828
rect 546552 3816 546558 3868
rect 273162 3748 273168 3800
rect 273220 3788 273226 3800
rect 293126 3788 293132 3800
rect 273220 3760 293132 3788
rect 273220 3748 273226 3760
rect 293126 3748 293132 3760
rect 293184 3748 293190 3800
rect 296622 3748 296628 3800
rect 296680 3788 296686 3800
rect 350258 3788 350264 3800
rect 296680 3760 350264 3788
rect 296680 3748 296686 3760
rect 350258 3748 350264 3760
rect 350316 3748 350322 3800
rect 376662 3748 376668 3800
rect 376720 3788 376726 3800
rect 550082 3788 550088 3800
rect 376720 3760 550088 3788
rect 376720 3748 376726 3760
rect 550082 3748 550088 3760
rect 550140 3748 550146 3800
rect 272996 3692 274220 3720
rect 34974 3612 34980 3664
rect 35032 3652 35038 3664
rect 36538 3652 36544 3664
rect 35032 3624 36544 3652
rect 35032 3612 35038 3624
rect 36538 3612 36544 3624
rect 36596 3612 36602 3664
rect 43346 3612 43352 3664
rect 43404 3652 43410 3664
rect 162121 3655 162179 3661
rect 162121 3652 162133 3655
rect 43404 3624 162133 3652
rect 43404 3612 43410 3624
rect 162121 3621 162133 3624
rect 162167 3621 162179 3655
rect 162121 3615 162179 3621
rect 162213 3655 162271 3661
rect 162213 3621 162225 3655
rect 162259 3652 162271 3655
rect 165798 3652 165804 3664
rect 162259 3624 165804 3652
rect 162259 3621 162271 3624
rect 162213 3615 162271 3621
rect 165798 3612 165804 3624
rect 165856 3612 165862 3664
rect 166997 3655 167055 3661
rect 166997 3621 167009 3655
rect 167043 3652 167055 3655
rect 170585 3655 170643 3661
rect 167043 3624 169892 3652
rect 167043 3621 167055 3624
rect 166997 3615 167055 3621
rect 39758 3544 39764 3596
rect 39816 3584 39822 3596
rect 169754 3584 169760 3596
rect 39816 3556 169760 3584
rect 39816 3544 39822 3556
rect 169754 3544 169760 3556
rect 169812 3544 169818 3596
rect 169864 3584 169892 3624
rect 170585 3621 170597 3655
rect 170631 3652 170643 3655
rect 182174 3652 182180 3664
rect 170631 3624 182180 3652
rect 170631 3621 170643 3624
rect 170585 3615 170643 3621
rect 182174 3612 182180 3624
rect 182232 3612 182238 3664
rect 193214 3612 193220 3664
rect 193272 3652 193278 3664
rect 194410 3652 194416 3664
rect 193272 3624 194416 3652
rect 193272 3612 193278 3624
rect 194410 3612 194416 3624
rect 194468 3612 194474 3664
rect 201405 3655 201463 3661
rect 201405 3621 201417 3655
rect 201451 3652 201463 3655
rect 202877 3655 202935 3661
rect 202877 3652 202889 3655
rect 201451 3624 202889 3652
rect 201451 3621 201463 3624
rect 201405 3615 201463 3621
rect 202877 3621 202889 3624
rect 202923 3621 202935 3655
rect 202877 3615 202935 3621
rect 207474 3612 207480 3664
rect 207532 3652 207538 3664
rect 237466 3652 237472 3664
rect 207532 3624 237472 3652
rect 207532 3612 207538 3624
rect 237466 3612 237472 3624
rect 237524 3612 237530 3664
rect 251358 3652 251364 3664
rect 249076 3624 251364 3652
rect 173989 3587 174047 3593
rect 173989 3584 174001 3587
rect 169864 3556 174001 3584
rect 173989 3553 174001 3556
rect 174035 3553 174047 3587
rect 173989 3547 174047 3553
rect 206097 3587 206155 3593
rect 206097 3553 206109 3587
rect 206143 3584 206155 3587
rect 226337 3587 226395 3593
rect 226337 3584 226349 3587
rect 206143 3556 226349 3584
rect 206143 3553 206155 3556
rect 206097 3547 206155 3553
rect 226337 3553 226349 3556
rect 226383 3553 226395 3587
rect 226337 3547 226395 3553
rect 226429 3587 226487 3593
rect 226429 3553 226441 3587
rect 226475 3584 226487 3587
rect 240410 3584 240416 3596
rect 226475 3556 240416 3584
rect 226475 3553 226487 3556
rect 226429 3547 226487 3553
rect 240410 3544 240416 3556
rect 240468 3544 240474 3596
rect 16022 3476 16028 3528
rect 16080 3516 16086 3528
rect 19978 3516 19984 3528
rect 16080 3488 19984 3516
rect 16080 3476 16086 3488
rect 19978 3476 19984 3488
rect 20036 3476 20042 3528
rect 25498 3476 25504 3528
rect 25556 3516 25562 3528
rect 29638 3516 29644 3528
rect 25556 3488 29644 3516
rect 25556 3476 25562 3488
rect 29638 3476 29644 3488
rect 29696 3476 29702 3528
rect 31478 3476 31484 3528
rect 31536 3516 31542 3528
rect 32398 3516 32404 3528
rect 31536 3488 32404 3516
rect 31536 3476 31542 3488
rect 32398 3476 32404 3488
rect 32456 3476 32462 3528
rect 32674 3476 32680 3528
rect 32732 3516 32738 3528
rect 35158 3516 35164 3528
rect 32732 3488 35164 3516
rect 32732 3476 32738 3488
rect 35158 3476 35164 3488
rect 35216 3476 35222 3528
rect 42150 3476 42156 3528
rect 42208 3516 42214 3528
rect 42702 3516 42708 3528
rect 42208 3488 42708 3516
rect 42208 3476 42214 3488
rect 42702 3476 42708 3488
rect 42760 3476 42766 3528
rect 42797 3519 42855 3525
rect 42797 3485 42809 3519
rect 42843 3516 42855 3519
rect 168742 3516 168748 3528
rect 42843 3488 168748 3516
rect 42843 3485 42855 3488
rect 42797 3479 42855 3485
rect 168742 3476 168748 3488
rect 168800 3476 168806 3528
rect 183738 3476 183744 3528
rect 183796 3516 183802 3528
rect 184842 3516 184848 3528
rect 183796 3488 184848 3516
rect 183796 3476 183802 3488
rect 184842 3476 184848 3488
rect 184900 3476 184906 3528
rect 202877 3519 202935 3525
rect 202877 3485 202889 3519
rect 202923 3516 202935 3519
rect 211157 3519 211215 3525
rect 211157 3516 211169 3519
rect 202923 3488 211169 3516
rect 202923 3485 202935 3488
rect 202877 3479 202935 3485
rect 211157 3485 211169 3488
rect 211203 3485 211215 3519
rect 211157 3479 211215 3485
rect 220725 3519 220783 3525
rect 220725 3485 220737 3519
rect 220771 3516 220783 3519
rect 230477 3519 230535 3525
rect 230477 3516 230489 3519
rect 220771 3488 230489 3516
rect 220771 3485 220783 3488
rect 220725 3479 220783 3485
rect 230477 3485 230489 3488
rect 230523 3485 230535 3519
rect 230477 3479 230535 3485
rect 233513 3519 233571 3525
rect 233513 3485 233525 3519
rect 233559 3516 233571 3519
rect 237558 3516 237564 3528
rect 233559 3488 237564 3516
rect 233559 3485 233571 3488
rect 233513 3479 233571 3485
rect 237558 3476 237564 3488
rect 237616 3476 237622 3528
rect 241974 3476 241980 3528
rect 242032 3516 242038 3528
rect 242802 3516 242808 3528
rect 242032 3488 242808 3516
rect 242032 3476 242038 3488
rect 242802 3476 242808 3488
rect 242860 3476 242866 3528
rect 249076 3516 249104 3624
rect 251358 3612 251364 3624
rect 251416 3612 251422 3664
rect 266170 3612 266176 3664
rect 266228 3652 266234 3664
rect 274082 3652 274088 3664
rect 266228 3624 274088 3652
rect 266228 3612 266234 3624
rect 274082 3612 274088 3624
rect 274140 3612 274146 3664
rect 274192 3652 274220 3692
rect 274542 3680 274548 3732
rect 274600 3720 274606 3732
rect 296714 3720 296720 3732
rect 274600 3692 296720 3720
rect 274600 3680 274606 3692
rect 296714 3680 296720 3692
rect 296772 3680 296778 3732
rect 298002 3680 298008 3732
rect 298060 3720 298066 3732
rect 298060 3692 300440 3720
rect 298060 3680 298066 3692
rect 275649 3655 275707 3661
rect 275649 3652 275661 3655
rect 274192 3624 275661 3652
rect 275649 3621 275661 3624
rect 275695 3621 275707 3655
rect 275649 3615 275707 3621
rect 275922 3612 275928 3664
rect 275980 3652 275986 3664
rect 300302 3652 300308 3664
rect 275980 3624 300308 3652
rect 275980 3612 275986 3624
rect 300302 3612 300308 3624
rect 300360 3612 300366 3664
rect 300412 3652 300440 3692
rect 300762 3680 300768 3732
rect 300820 3720 300826 3732
rect 300820 3692 304948 3720
rect 300820 3680 300826 3692
rect 304813 3655 304871 3661
rect 304813 3652 304825 3655
rect 300412 3624 304825 3652
rect 304813 3621 304825 3624
rect 304859 3621 304871 3655
rect 304920 3652 304948 3692
rect 304994 3680 305000 3732
rect 305052 3720 305058 3732
rect 306098 3720 306104 3732
rect 305052 3692 306104 3720
rect 305052 3680 305058 3692
rect 306098 3680 306104 3692
rect 306156 3680 306162 3732
rect 306285 3723 306343 3729
rect 306285 3689 306297 3723
rect 306331 3720 306343 3723
rect 353754 3720 353760 3732
rect 306331 3692 353760 3720
rect 306331 3689 306343 3692
rect 306285 3683 306343 3689
rect 353754 3680 353760 3692
rect 353812 3680 353818 3732
rect 378042 3680 378048 3732
rect 378100 3720 378106 3732
rect 553578 3720 553584 3732
rect 378100 3692 553584 3720
rect 378100 3680 378106 3692
rect 553578 3680 553584 3692
rect 553636 3680 553642 3732
rect 360930 3652 360936 3664
rect 304920 3624 360936 3652
rect 304813 3615 304871 3621
rect 360930 3612 360936 3624
rect 360988 3612 360994 3664
rect 379422 3612 379428 3664
rect 379480 3652 379486 3664
rect 557166 3652 557172 3664
rect 379480 3624 557172 3652
rect 379480 3612 379486 3624
rect 557166 3612 557172 3624
rect 557224 3612 557230 3664
rect 266262 3544 266268 3596
rect 266320 3584 266326 3596
rect 276474 3584 276480 3596
rect 266320 3556 276480 3584
rect 266320 3544 266326 3556
rect 276474 3544 276480 3556
rect 276532 3544 276538 3596
rect 277302 3544 277308 3596
rect 277360 3584 277366 3596
rect 303798 3584 303804 3596
rect 277360 3556 303804 3584
rect 277360 3544 277366 3556
rect 303798 3544 303804 3556
rect 303856 3544 303862 3596
rect 304902 3544 304908 3596
rect 304960 3584 304966 3596
rect 306101 3587 306159 3593
rect 306101 3584 306113 3587
rect 304960 3556 306113 3584
rect 304960 3544 304966 3556
rect 306101 3553 306113 3556
rect 306147 3553 306159 3587
rect 306101 3547 306159 3553
rect 306285 3587 306343 3593
rect 306285 3553 306297 3587
rect 306331 3584 306343 3587
rect 371602 3584 371608 3596
rect 306331 3556 371608 3584
rect 306331 3553 306343 3556
rect 306285 3547 306343 3553
rect 371602 3544 371608 3556
rect 371660 3544 371666 3596
rect 380802 3544 380808 3596
rect 380860 3584 380866 3596
rect 560754 3584 560760 3596
rect 380860 3556 560760 3584
rect 380860 3544 380866 3556
rect 560754 3544 560760 3556
rect 560812 3544 560818 3596
rect 242912 3488 249104 3516
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 10318 3448 10324 3460
rect 6512 3420 10324 3448
rect 6512 3408 6518 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 29086 3408 29092 3460
rect 29144 3448 29150 3460
rect 162029 3451 162087 3457
rect 162029 3448 162041 3451
rect 29144 3420 162041 3448
rect 29144 3408 29150 3420
rect 162029 3417 162041 3420
rect 162075 3417 162087 3451
rect 162029 3411 162087 3417
rect 162121 3451 162179 3457
rect 162121 3417 162133 3451
rect 162167 3448 162179 3451
rect 171134 3448 171140 3460
rect 162167 3420 171140 3448
rect 162167 3417 162179 3420
rect 162121 3411 162179 3417
rect 171134 3408 171140 3420
rect 171192 3408 171198 3460
rect 189626 3408 189632 3460
rect 189684 3448 189690 3460
rect 189684 3420 205496 3448
rect 189684 3408 189690 3420
rect 45738 3340 45744 3392
rect 45796 3380 45802 3392
rect 46842 3380 46848 3392
rect 45796 3352 46848 3380
rect 45796 3340 45802 3352
rect 46842 3340 46848 3352
rect 46900 3340 46906 3392
rect 50522 3340 50528 3392
rect 50580 3380 50586 3392
rect 50982 3380 50988 3392
rect 50580 3352 50988 3380
rect 50580 3340 50586 3352
rect 50982 3340 50988 3352
rect 51040 3340 51046 3392
rect 54018 3340 54024 3392
rect 54076 3380 54082 3392
rect 55122 3380 55128 3392
rect 54076 3352 55128 3380
rect 54076 3340 54082 3352
rect 55122 3340 55128 3352
rect 55180 3340 55186 3392
rect 61194 3340 61200 3392
rect 61252 3380 61258 3392
rect 62022 3380 62028 3392
rect 61252 3352 62028 3380
rect 61252 3340 61258 3352
rect 62022 3340 62028 3352
rect 62080 3340 62086 3392
rect 81434 3340 81440 3392
rect 81492 3380 81498 3392
rect 82722 3380 82728 3392
rect 81492 3352 82728 3380
rect 81492 3340 81498 3352
rect 82722 3340 82728 3352
rect 82780 3340 82786 3392
rect 84841 3383 84899 3389
rect 84841 3380 84853 3383
rect 82832 3352 84853 3380
rect 18322 3272 18328 3324
rect 18380 3312 18386 3324
rect 21358 3312 21364 3324
rect 18380 3284 21364 3312
rect 18380 3272 18386 3284
rect 21358 3272 21364 3284
rect 21416 3272 21422 3324
rect 36170 3272 36176 3324
rect 36228 3312 36234 3324
rect 42797 3315 42855 3321
rect 42797 3312 42809 3315
rect 36228 3284 42809 3312
rect 36228 3272 36234 3284
rect 42797 3281 42809 3284
rect 42843 3281 42855 3315
rect 42797 3275 42855 3281
rect 27890 3204 27896 3256
rect 27948 3244 27954 3256
rect 31018 3244 31024 3256
rect 27948 3216 31024 3244
rect 27948 3204 27954 3216
rect 31018 3204 31024 3216
rect 31076 3204 31082 3256
rect 79042 3204 79048 3256
rect 79100 3244 79106 3256
rect 82832 3244 82860 3352
rect 84841 3349 84853 3352
rect 84887 3349 84899 3383
rect 84841 3343 84899 3349
rect 84930 3340 84936 3392
rect 84988 3380 84994 3392
rect 85482 3380 85488 3392
rect 84988 3352 85488 3380
rect 84988 3340 84994 3352
rect 85482 3340 85488 3352
rect 85540 3340 85546 3392
rect 88518 3340 88524 3392
rect 88576 3380 88582 3392
rect 89622 3380 89628 3392
rect 88576 3352 89628 3380
rect 88576 3340 88582 3352
rect 89622 3340 89628 3352
rect 89680 3340 89686 3392
rect 189074 3380 189080 3392
rect 89824 3352 189080 3380
rect 79100 3216 82860 3244
rect 79100 3204 79106 3216
rect 86126 3204 86132 3256
rect 86184 3244 86190 3256
rect 89824 3244 89852 3352
rect 189074 3340 189080 3352
rect 189132 3340 189138 3392
rect 205468 3380 205496 3420
rect 212258 3408 212264 3460
rect 212316 3448 212322 3460
rect 224865 3451 224923 3457
rect 224865 3448 224877 3451
rect 212316 3420 224877 3448
rect 212316 3408 212322 3420
rect 224865 3417 224877 3420
rect 224911 3417 224923 3451
rect 224865 3411 224923 3417
rect 239582 3408 239588 3460
rect 239640 3448 239646 3460
rect 242912 3448 242940 3488
rect 249150 3476 249156 3528
rect 249208 3516 249214 3528
rect 249702 3516 249708 3528
rect 249208 3488 249708 3516
rect 249208 3476 249214 3488
rect 249702 3476 249708 3488
rect 249760 3476 249766 3528
rect 252646 3476 252652 3528
rect 252704 3516 252710 3528
rect 253842 3516 253848 3528
rect 252704 3488 253848 3516
rect 252704 3476 252710 3488
rect 253842 3476 253848 3488
rect 253900 3476 253906 3528
rect 267642 3476 267648 3528
rect 267700 3516 267706 3528
rect 277670 3516 277676 3528
rect 267700 3488 277676 3516
rect 267700 3476 267706 3488
rect 277670 3476 277676 3488
rect 277728 3476 277734 3528
rect 280062 3476 280068 3528
rect 280120 3516 280126 3528
rect 307386 3516 307392 3528
rect 280120 3488 307392 3516
rect 280120 3476 280126 3488
rect 307386 3476 307392 3488
rect 307444 3476 307450 3528
rect 309042 3476 309048 3528
rect 309100 3516 309106 3528
rect 382366 3516 382372 3528
rect 309100 3488 382372 3516
rect 309100 3476 309106 3488
rect 382366 3476 382372 3488
rect 382424 3476 382430 3528
rect 384942 3476 384948 3528
rect 385000 3516 385006 3528
rect 567838 3516 567844 3528
rect 385000 3488 567844 3516
rect 385000 3476 385006 3488
rect 567838 3476 567844 3488
rect 567896 3476 567902 3528
rect 239640 3420 242940 3448
rect 242989 3451 243047 3457
rect 239640 3408 239646 3420
rect 242989 3417 243001 3451
rect 243035 3448 243047 3451
rect 249886 3448 249892 3460
rect 243035 3420 249892 3448
rect 243035 3417 243047 3420
rect 242989 3411 243047 3417
rect 249886 3408 249892 3420
rect 249944 3408 249950 3460
rect 267550 3408 267556 3460
rect 267608 3448 267614 3460
rect 278866 3448 278872 3460
rect 267608 3420 278872 3448
rect 267608 3408 267614 3420
rect 278866 3408 278872 3420
rect 278924 3408 278930 3460
rect 281442 3408 281448 3460
rect 281500 3448 281506 3460
rect 310974 3448 310980 3460
rect 281500 3420 310980 3448
rect 281500 3408 281506 3420
rect 310974 3408 310980 3420
rect 311032 3408 311038 3460
rect 311802 3408 311808 3460
rect 311860 3448 311866 3460
rect 389450 3448 389456 3460
rect 311860 3420 389456 3448
rect 311860 3408 311866 3420
rect 389450 3408 389456 3420
rect 389508 3408 389514 3460
rect 390462 3408 390468 3460
rect 390520 3448 390526 3460
rect 582190 3448 582196 3460
rect 390520 3420 582196 3448
rect 390520 3408 390526 3420
rect 582190 3408 582196 3420
rect 582248 3408 582254 3460
rect 205468 3352 205680 3380
rect 89898 3272 89904 3324
rect 89956 3312 89962 3324
rect 190730 3312 190736 3324
rect 89956 3284 190736 3312
rect 89956 3272 89962 3284
rect 190730 3272 190736 3284
rect 190788 3272 190794 3324
rect 205652 3312 205680 3352
rect 225322 3340 225328 3392
rect 225380 3380 225386 3392
rect 245746 3380 245752 3392
rect 225380 3352 245752 3380
rect 225380 3340 225386 3352
rect 245746 3340 245752 3352
rect 245804 3340 245810 3392
rect 269022 3340 269028 3392
rect 269080 3380 269086 3392
rect 275649 3383 275707 3389
rect 269080 3352 275416 3380
rect 269080 3340 269086 3352
rect 205652 3284 215340 3312
rect 86184 3216 89852 3244
rect 86184 3204 86190 3216
rect 93302 3204 93308 3256
rect 93360 3244 93366 3256
rect 192110 3244 192116 3256
rect 93360 3216 192116 3244
rect 93360 3204 93366 3216
rect 192110 3204 192116 3216
rect 192168 3204 192174 3256
rect 84749 3179 84807 3185
rect 84749 3145 84761 3179
rect 84795 3176 84807 3179
rect 93765 3179 93823 3185
rect 93765 3176 93777 3179
rect 84795 3148 93777 3176
rect 84795 3145 84807 3148
rect 84749 3139 84807 3145
rect 93765 3145 93777 3148
rect 93811 3145 93823 3179
rect 93765 3139 93823 3145
rect 95694 3136 95700 3188
rect 95752 3176 95758 3188
rect 96522 3176 96528 3188
rect 95752 3148 96528 3176
rect 95752 3136 95758 3148
rect 96522 3136 96528 3148
rect 96580 3136 96586 3188
rect 102778 3136 102784 3188
rect 102836 3176 102842 3188
rect 103422 3176 103428 3188
rect 102836 3148 103428 3176
rect 102836 3136 102842 3148
rect 103422 3136 103428 3148
rect 103480 3136 103486 3188
rect 106366 3136 106372 3188
rect 106424 3176 106430 3188
rect 107562 3176 107568 3188
rect 106424 3148 107568 3176
rect 106424 3136 106430 3148
rect 107562 3136 107568 3148
rect 107620 3136 107626 3188
rect 107657 3179 107715 3185
rect 107657 3145 107669 3179
rect 107703 3176 107715 3179
rect 111061 3179 111119 3185
rect 111061 3176 111073 3179
rect 107703 3148 111073 3176
rect 107703 3145 107715 3148
rect 107657 3139 107715 3145
rect 111061 3145 111073 3148
rect 111107 3145 111119 3179
rect 111061 3139 111119 3145
rect 111150 3136 111156 3188
rect 111208 3176 111214 3188
rect 111702 3176 111708 3188
rect 111208 3148 111708 3176
rect 111208 3136 111214 3148
rect 111702 3136 111708 3148
rect 111760 3136 111766 3188
rect 111797 3179 111855 3185
rect 111797 3145 111809 3179
rect 111843 3176 111855 3179
rect 193398 3176 193404 3188
rect 111843 3148 193404 3176
rect 111843 3145 111855 3148
rect 111797 3139 111855 3145
rect 193398 3136 193404 3148
rect 193456 3136 193462 3188
rect 100478 3068 100484 3120
rect 100536 3108 100542 3120
rect 194594 3108 194600 3120
rect 100536 3080 194600 3108
rect 100536 3068 100542 3080
rect 194594 3068 194600 3080
rect 194652 3068 194658 3120
rect 96890 3000 96896 3052
rect 96948 3040 96954 3052
rect 111797 3043 111855 3049
rect 111797 3040 111809 3043
rect 96948 3012 111809 3040
rect 96948 3000 96954 3012
rect 111797 3009 111809 3012
rect 111843 3009 111855 3043
rect 111797 3003 111855 3009
rect 111889 3043 111947 3049
rect 111889 3009 111901 3043
rect 111935 3040 111947 3043
rect 196158 3040 196164 3052
rect 111935 3012 196164 3040
rect 111935 3009 111947 3012
rect 111889 3003 111947 3009
rect 196158 3000 196164 3012
rect 196216 3000 196222 3052
rect 196802 3000 196808 3052
rect 196860 3040 196866 3052
rect 197262 3040 197268 3052
rect 196860 3012 197268 3040
rect 196860 3000 196866 3012
rect 197262 3000 197268 3012
rect 197320 3000 197326 3052
rect 215312 3040 215340 3284
rect 227714 3272 227720 3324
rect 227772 3312 227778 3324
rect 229002 3312 229008 3324
rect 227772 3284 229008 3312
rect 227772 3272 227778 3284
rect 229002 3272 229008 3284
rect 229060 3272 229066 3324
rect 247126 3312 247132 3324
rect 229112 3284 247132 3312
rect 228910 3204 228916 3256
rect 228968 3244 228974 3256
rect 229112 3244 229140 3284
rect 247126 3272 247132 3284
rect 247184 3272 247190 3324
rect 268378 3272 268384 3324
rect 268436 3312 268442 3324
rect 275278 3312 275284 3324
rect 268436 3284 275284 3312
rect 268436 3272 268442 3284
rect 275278 3272 275284 3284
rect 275336 3272 275342 3324
rect 275388 3312 275416 3352
rect 275649 3349 275661 3383
rect 275695 3380 275707 3383
rect 282454 3380 282460 3392
rect 275695 3352 282460 3380
rect 275695 3349 275707 3352
rect 275649 3343 275707 3349
rect 282454 3340 282460 3352
rect 282512 3340 282518 3392
rect 286870 3340 286876 3392
rect 286928 3380 286934 3392
rect 327626 3380 327632 3392
rect 286928 3352 327632 3380
rect 286928 3340 286934 3352
rect 327626 3340 327632 3352
rect 327684 3340 327690 3392
rect 336642 3340 336648 3392
rect 336700 3380 336706 3392
rect 450170 3380 450176 3392
rect 336700 3352 450176 3380
rect 336700 3340 336706 3352
rect 450170 3340 450176 3352
rect 450228 3340 450234 3392
rect 459554 3340 459560 3392
rect 459612 3380 459618 3392
rect 460842 3380 460848 3392
rect 459612 3352 460848 3380
rect 459612 3340 459618 3352
rect 460842 3340 460848 3352
rect 460900 3340 460906 3392
rect 281258 3312 281264 3324
rect 275388 3284 281264 3312
rect 281258 3272 281264 3284
rect 281316 3272 281322 3324
rect 288158 3272 288164 3324
rect 288216 3312 288222 3324
rect 328822 3312 328828 3324
rect 288216 3284 328828 3312
rect 288216 3272 288222 3284
rect 328822 3272 328828 3284
rect 328880 3272 328886 3324
rect 333882 3272 333888 3324
rect 333940 3312 333946 3324
rect 442994 3312 443000 3324
rect 333940 3284 443000 3312
rect 333940 3272 333946 3284
rect 442994 3272 443000 3284
rect 443052 3272 443058 3324
rect 228968 3216 229140 3244
rect 228968 3204 228974 3216
rect 232498 3204 232504 3256
rect 232556 3244 232562 3256
rect 232556 3216 234660 3244
rect 232556 3204 232562 3216
rect 224126 3136 224132 3188
rect 224184 3176 224190 3188
rect 232406 3176 232412 3188
rect 224184 3148 232412 3176
rect 224184 3136 224190 3148
rect 232406 3136 232412 3148
rect 232464 3136 232470 3188
rect 234632 3108 234660 3216
rect 235994 3204 236000 3256
rect 236052 3244 236058 3256
rect 242989 3247 243047 3253
rect 242989 3244 243001 3247
rect 236052 3216 243001 3244
rect 236052 3204 236058 3216
rect 242989 3213 243001 3216
rect 243035 3213 243047 3247
rect 242989 3207 243047 3213
rect 251450 3204 251456 3256
rect 251508 3244 251514 3256
rect 254578 3244 254584 3256
rect 251508 3216 254584 3244
rect 251508 3204 251514 3216
rect 254578 3204 254584 3216
rect 254636 3204 254642 3256
rect 280062 3244 280068 3256
rect 275572 3216 280068 3244
rect 253842 3136 253848 3188
rect 253900 3176 253906 3188
rect 257062 3176 257068 3188
rect 253900 3148 257068 3176
rect 253900 3136 253906 3148
rect 257062 3136 257068 3148
rect 257120 3136 257126 3188
rect 243538 3108 243544 3120
rect 234632 3080 243544 3108
rect 243538 3068 243544 3080
rect 243596 3068 243602 3120
rect 250346 3068 250352 3120
rect 250404 3108 250410 3120
rect 251082 3108 251088 3120
rect 250404 3080 251088 3108
rect 250404 3068 250410 3080
rect 251082 3068 251088 3080
rect 251140 3068 251146 3120
rect 268930 3068 268936 3120
rect 268988 3108 268994 3120
rect 275572 3108 275600 3216
rect 280062 3204 280068 3216
rect 280120 3204 280126 3256
rect 285582 3204 285588 3256
rect 285640 3244 285646 3256
rect 285640 3216 320036 3244
rect 285640 3204 285646 3216
rect 286962 3136 286968 3188
rect 287020 3176 287026 3188
rect 319901 3179 319959 3185
rect 319901 3176 319913 3179
rect 287020 3148 319913 3176
rect 287020 3136 287026 3148
rect 319901 3145 319913 3148
rect 319947 3145 319959 3179
rect 320008 3176 320036 3216
rect 321646 3204 321652 3256
rect 321704 3244 321710 3256
rect 322842 3244 322848 3256
rect 321704 3216 322848 3244
rect 321704 3204 321710 3216
rect 322842 3204 322848 3216
rect 322900 3204 322906 3256
rect 331122 3204 331128 3256
rect 331180 3244 331186 3256
rect 435818 3244 435824 3256
rect 331180 3216 435824 3244
rect 331180 3204 331186 3216
rect 435818 3204 435824 3216
rect 435876 3204 435882 3256
rect 324038 3176 324044 3188
rect 320008 3148 324044 3176
rect 319901 3139 319959 3145
rect 324038 3136 324044 3148
rect 324096 3136 324102 3188
rect 328362 3136 328368 3188
rect 328420 3176 328426 3188
rect 428734 3176 428740 3188
rect 328420 3148 428740 3176
rect 328420 3136 328426 3148
rect 428734 3136 428740 3148
rect 428792 3136 428798 3188
rect 268988 3080 275600 3108
rect 268988 3068 268994 3080
rect 285490 3068 285496 3120
rect 285548 3108 285554 3120
rect 321646 3108 321652 3120
rect 285548 3080 321652 3108
rect 285548 3068 285554 3080
rect 321646 3068 321652 3080
rect 321704 3068 321710 3120
rect 325421 3111 325479 3117
rect 325421 3108 325433 3111
rect 321756 3080 325433 3108
rect 222197 3043 222255 3049
rect 222197 3040 222209 3043
rect 215312 3012 222209 3040
rect 222197 3009 222209 3012
rect 222243 3009 222255 3043
rect 222197 3003 222255 3009
rect 226337 3043 226395 3049
rect 226337 3009 226349 3043
rect 226383 3040 226395 3043
rect 233513 3043 233571 3049
rect 233513 3040 233525 3043
rect 226383 3012 233525 3040
rect 226383 3009 226395 3012
rect 226337 3003 226395 3009
rect 233513 3009 233525 3012
rect 233559 3009 233571 3043
rect 233513 3003 233571 3009
rect 262858 3000 262864 3052
rect 262916 3040 262922 3052
rect 264606 3040 264612 3052
rect 262916 3012 264612 3040
rect 262916 3000 262922 3012
rect 264606 3000 264612 3012
rect 264664 3000 264670 3052
rect 284110 3000 284116 3052
rect 284168 3040 284174 3052
rect 320450 3040 320456 3052
rect 284168 3012 320456 3040
rect 284168 3000 284174 3012
rect 320450 3000 320456 3012
rect 320508 3000 320514 3052
rect 320545 3043 320603 3049
rect 320545 3009 320557 3043
rect 320591 3040 320603 3043
rect 321756 3040 321784 3080
rect 325421 3077 325433 3080
rect 325467 3077 325479 3111
rect 325421 3071 325479 3077
rect 325602 3068 325608 3120
rect 325660 3108 325666 3120
rect 325660 3080 416728 3108
rect 325660 3068 325666 3080
rect 320591 3012 321784 3040
rect 320591 3009 320603 3012
rect 320545 3003 320603 3009
rect 322750 3000 322756 3052
rect 322808 3040 322814 3052
rect 414474 3040 414480 3052
rect 322808 3012 414480 3040
rect 322808 3000 322814 3012
rect 414474 3000 414480 3012
rect 414532 3000 414538 3052
rect 416700 3040 416728 3080
rect 416774 3068 416780 3120
rect 416832 3108 416838 3120
rect 417970 3108 417976 3120
rect 416832 3080 417976 3108
rect 416832 3068 416838 3080
rect 417970 3068 417976 3080
rect 418028 3068 418034 3120
rect 421558 3040 421564 3052
rect 416700 3012 421564 3040
rect 421558 3000 421564 3012
rect 421616 3000 421622 3052
rect 10042 2932 10048 2984
rect 10100 2972 10106 2984
rect 11698 2972 11704 2984
rect 10100 2944 11704 2972
rect 10100 2932 10106 2944
rect 11698 2932 11704 2944
rect 11756 2932 11762 2984
rect 24302 2932 24308 2984
rect 24360 2972 24366 2984
rect 28258 2972 28264 2984
rect 24360 2944 28264 2972
rect 24360 2932 24366 2944
rect 28258 2932 28264 2944
rect 28316 2932 28322 2984
rect 113542 2932 113548 2984
rect 113600 2972 113606 2984
rect 114462 2972 114468 2984
rect 113600 2944 114468 2972
rect 113600 2932 113606 2944
rect 114462 2932 114468 2944
rect 114520 2932 114526 2984
rect 120626 2932 120632 2984
rect 120684 2972 120690 2984
rect 121362 2972 121368 2984
rect 120684 2944 121368 2972
rect 120684 2932 120690 2944
rect 121362 2932 121368 2944
rect 121420 2932 121426 2984
rect 197630 2972 197636 2984
rect 121564 2944 197636 2972
rect 114738 2864 114744 2916
rect 114796 2904 114802 2916
rect 121457 2907 121515 2913
rect 121457 2904 121469 2907
rect 114796 2876 121469 2904
rect 114796 2864 114802 2876
rect 121457 2873 121469 2876
rect 121503 2873 121515 2907
rect 121457 2867 121515 2873
rect 103974 2796 103980 2848
rect 104032 2836 104038 2848
rect 107473 2839 107531 2845
rect 107473 2836 107485 2839
rect 104032 2808 107485 2836
rect 104032 2796 104038 2808
rect 107473 2805 107485 2808
rect 107519 2805 107531 2839
rect 107473 2799 107531 2805
rect 107562 2796 107568 2848
rect 107620 2836 107626 2848
rect 121564 2836 121592 2944
rect 197630 2932 197636 2944
rect 197688 2932 197694 2984
rect 231302 2932 231308 2984
rect 231360 2972 231366 2984
rect 235258 2972 235264 2984
rect 231360 2944 235264 2972
rect 231360 2932 231366 2944
rect 235258 2932 235264 2944
rect 235316 2932 235322 2984
rect 263502 2932 263508 2984
rect 263560 2972 263566 2984
rect 269298 2972 269304 2984
rect 263560 2944 269304 2972
rect 263560 2932 263566 2944
rect 269298 2932 269304 2944
rect 269356 2932 269362 2984
rect 282730 2932 282736 2984
rect 282788 2972 282794 2984
rect 316954 2972 316960 2984
rect 282788 2944 316960 2972
rect 282788 2932 282794 2944
rect 316954 2932 316960 2944
rect 317012 2932 317018 2984
rect 317322 2932 317328 2984
rect 317380 2972 317386 2984
rect 319901 2975 319959 2981
rect 317380 2944 318196 2972
rect 317380 2932 317386 2944
rect 121641 2907 121699 2913
rect 121641 2873 121653 2907
rect 121687 2904 121699 2907
rect 200298 2904 200304 2916
rect 121687 2876 200304 2904
rect 121687 2873 121699 2876
rect 121641 2867 121699 2873
rect 200298 2864 200304 2876
rect 200356 2864 200362 2916
rect 245562 2864 245568 2916
rect 245620 2904 245626 2916
rect 246298 2904 246304 2916
rect 245620 2876 246304 2904
rect 245620 2864 245626 2876
rect 246298 2864 246304 2876
rect 246356 2864 246362 2916
rect 284202 2864 284208 2916
rect 284260 2904 284266 2916
rect 318058 2904 318064 2916
rect 284260 2876 318064 2904
rect 284260 2864 284266 2876
rect 318058 2864 318064 2876
rect 318116 2864 318122 2916
rect 318168 2904 318196 2944
rect 319901 2941 319913 2975
rect 319947 2972 319959 2975
rect 325234 2972 325240 2984
rect 319947 2944 325240 2972
rect 319947 2941 319959 2944
rect 319901 2935 319959 2941
rect 325234 2932 325240 2944
rect 325292 2932 325298 2984
rect 407298 2972 407304 2984
rect 325344 2944 407304 2972
rect 319993 2907 320051 2913
rect 319993 2904 320005 2907
rect 318168 2876 320005 2904
rect 319993 2873 320005 2876
rect 320039 2873 320051 2907
rect 319993 2867 320051 2873
rect 320082 2864 320088 2916
rect 320140 2904 320146 2916
rect 325344 2904 325372 2944
rect 407298 2932 407304 2944
rect 407356 2932 407362 2984
rect 320140 2876 325372 2904
rect 325421 2907 325479 2913
rect 320140 2864 320146 2876
rect 325421 2873 325433 2907
rect 325467 2904 325479 2907
rect 400214 2904 400220 2916
rect 325467 2876 400220 2904
rect 325467 2873 325479 2876
rect 325421 2867 325479 2873
rect 400214 2864 400220 2876
rect 400272 2864 400278 2916
rect 107620 2808 121592 2836
rect 107620 2796 107626 2808
rect 121822 2796 121828 2848
rect 121880 2836 121886 2848
rect 122742 2836 122748 2848
rect 121880 2808 122748 2836
rect 121880 2796 121886 2808
rect 122742 2796 122748 2808
rect 122800 2796 122806 2848
rect 124214 2796 124220 2848
rect 124272 2836 124278 2848
rect 125502 2836 125508 2848
rect 124272 2808 125508 2836
rect 124272 2796 124278 2808
rect 125502 2796 125508 2808
rect 125560 2796 125566 2848
rect 125612 2808 127756 2836
rect 125410 2728 125416 2780
rect 125468 2768 125474 2780
rect 125612 2768 125640 2808
rect 125468 2740 125640 2768
rect 127728 2768 127756 2808
rect 127802 2796 127808 2848
rect 127860 2836 127866 2848
rect 128262 2836 128268 2848
rect 127860 2808 128268 2836
rect 127860 2796 127866 2808
rect 128262 2796 128268 2808
rect 128320 2796 128326 2848
rect 128372 2808 130148 2836
rect 128372 2768 128400 2808
rect 127728 2740 128400 2768
rect 130120 2768 130148 2808
rect 130194 2796 130200 2848
rect 130252 2836 130258 2848
rect 131022 2836 131028 2848
rect 130252 2808 131028 2836
rect 130252 2796 130258 2808
rect 131022 2796 131028 2808
rect 131080 2796 131086 2848
rect 131390 2796 131396 2848
rect 131448 2836 131454 2848
rect 132310 2836 132316 2848
rect 131448 2808 132316 2836
rect 131448 2796 131454 2808
rect 132310 2796 132316 2808
rect 132368 2796 132374 2848
rect 204254 2836 204260 2848
rect 132420 2808 204260 2836
rect 132420 2768 132448 2808
rect 204254 2796 204260 2808
rect 204312 2796 204318 2848
rect 255041 2839 255099 2845
rect 255041 2805 255053 2839
rect 255087 2836 255099 2839
rect 255222 2836 255228 2848
rect 255087 2808 255228 2836
rect 255087 2805 255099 2808
rect 255041 2799 255099 2805
rect 255222 2796 255228 2808
rect 255280 2796 255286 2848
rect 256234 2796 256240 2848
rect 256292 2836 256298 2848
rect 256602 2836 256608 2848
rect 256292 2808 256608 2836
rect 256292 2796 256298 2808
rect 256602 2796 256608 2808
rect 256660 2796 256666 2848
rect 282822 2796 282828 2848
rect 282880 2836 282886 2848
rect 314562 2836 314568 2848
rect 282880 2808 314568 2836
rect 282880 2796 282886 2808
rect 314562 2796 314568 2808
rect 314620 2796 314626 2848
rect 314654 2796 314660 2848
rect 314712 2836 314718 2848
rect 393038 2836 393044 2848
rect 314712 2808 393044 2836
rect 314712 2796 314718 2808
rect 393038 2796 393044 2808
rect 393096 2796 393102 2848
rect 130120 2740 132448 2768
rect 125468 2728 125474 2740
rect 385126 2592 385132 2644
rect 385184 2632 385190 2644
rect 385862 2632 385868 2644
rect 385184 2604 385868 2632
rect 385184 2592 385190 2604
rect 385862 2592 385868 2604
rect 385920 2592 385926 2644
rect 195606 1844 195612 1896
rect 195664 1884 195670 1896
rect 201405 1887 201463 1893
rect 201405 1884 201417 1887
rect 195664 1856 201417 1884
rect 195664 1844 195670 1856
rect 201405 1853 201417 1856
rect 201451 1853 201463 1887
rect 201405 1847 201463 1853
rect 205082 1232 205088 1284
rect 205140 1272 205146 1284
rect 206097 1275 206155 1281
rect 206097 1272 206109 1275
rect 205140 1244 206109 1272
rect 205140 1232 205146 1244
rect 206097 1241 206109 1244
rect 206143 1241 206155 1275
rect 206097 1235 206155 1241
rect 137278 552 137284 604
rect 137336 592 137342 604
rect 137922 592 137928 604
rect 137336 564 137928 592
rect 137336 552 137342 564
rect 137922 552 137928 564
rect 137980 552 137986 604
rect 138474 552 138480 604
rect 138532 592 138538 604
rect 139302 592 139308 604
rect 138532 564 139308 592
rect 138532 552 138538 564
rect 139302 552 139308 564
rect 139360 552 139366 604
rect 145650 552 145656 604
rect 145708 592 145714 604
rect 146202 592 146208 604
rect 145708 564 146208 592
rect 145708 552 145714 564
rect 146202 552 146208 564
rect 146260 552 146266 604
rect 148042 552 148048 604
rect 148100 592 148106 604
rect 148962 592 148968 604
rect 148100 564 148968 592
rect 148100 552 148106 564
rect 148962 552 148968 564
rect 149020 552 149026 604
rect 149238 552 149244 604
rect 149296 592 149302 604
rect 150342 592 150348 604
rect 149296 564 150348 592
rect 149296 552 149302 564
rect 150342 552 150348 564
rect 150400 552 150406 604
rect 151538 552 151544 604
rect 151596 592 151602 604
rect 151722 592 151728 604
rect 151596 564 151728 592
rect 151596 552 151602 564
rect 151722 552 151728 564
rect 151780 552 151786 604
rect 156322 552 156328 604
rect 156380 592 156386 604
rect 157242 592 157248 604
rect 156380 564 157248 592
rect 156380 552 156386 564
rect 157242 552 157248 564
rect 157300 552 157306 604
rect 187234 552 187240 604
rect 187292 592 187298 604
rect 187602 592 187608 604
rect 187292 564 187608 592
rect 187292 552 187298 564
rect 187602 552 187608 564
rect 187660 552 187666 604
rect 255038 592 255044 604
rect 254999 564 255044 592
rect 255038 552 255044 564
rect 255096 552 255102 604
rect 259638 552 259644 604
rect 259696 592 259702 604
rect 259822 592 259828 604
rect 259696 564 259828 592
rect 259696 552 259702 564
rect 259822 552 259828 564
rect 259880 552 259886 604
rect 265250 552 265256 604
rect 265308 592 265314 604
rect 265802 592 265808 604
rect 265308 564 265808 592
rect 265308 552 265314 564
rect 265802 552 265808 564
rect 265860 552 265866 604
rect 300854 552 300860 604
rect 300912 592 300918 604
rect 301406 592 301412 604
rect 300912 564 301412 592
rect 300912 552 300918 564
rect 301406 552 301412 564
rect 301464 552 301470 604
rect 307754 552 307760 604
rect 307812 592 307818 604
rect 308582 592 308588 604
rect 307812 564 308588 592
rect 307812 552 307818 564
rect 308582 552 308588 564
rect 308640 552 308646 604
rect 309134 552 309140 604
rect 309192 592 309198 604
rect 309778 592 309784 604
rect 309192 564 309784 592
rect 309192 552 309198 564
rect 309778 552 309784 564
rect 309836 552 309842 604
rect 314746 552 314752 604
rect 314804 592 314810 604
rect 315758 592 315764 604
rect 314804 564 315764 592
rect 314804 552 314810 564
rect 315758 552 315764 564
rect 315816 552 315822 604
rect 325694 552 325700 604
rect 325752 592 325758 604
rect 326430 592 326436 604
rect 325752 564 326436 592
rect 325752 552 325758 564
rect 326430 552 326436 564
rect 326488 552 326494 604
rect 332594 552 332600 604
rect 332652 592 332658 604
rect 333606 592 333612 604
rect 332652 564 333612 592
rect 332652 552 332658 564
rect 333606 552 333612 564
rect 333664 552 333670 604
rect 336734 552 336740 604
rect 336792 592 336798 604
rect 337102 592 337108 604
rect 336792 564 337108 592
rect 336792 552 336798 564
rect 337102 552 337108 564
rect 337160 552 337166 604
rect 339586 552 339592 604
rect 339644 592 339650 604
rect 340690 592 340696 604
rect 339644 564 340696 592
rect 339644 552 339650 564
rect 340690 552 340696 564
rect 340748 552 340754 604
rect 378134 552 378140 604
rect 378192 592 378198 604
rect 378778 592 378784 604
rect 378192 564 378784 592
rect 378192 552 378198 564
rect 378778 552 378784 564
rect 378836 552 378842 604
rect 520366 552 520372 604
rect 520424 592 520430 604
rect 521470 592 521476 604
rect 520424 564 521476 592
rect 520424 552 520430 564
rect 521470 552 521476 564
rect 521528 552 521534 604
rect 524414 552 524420 604
rect 524472 592 524478 604
rect 525058 592 525064 604
rect 524472 564 525064 592
rect 524472 552 524478 564
rect 525058 552 525064 564
rect 525116 552 525122 604
rect 531314 552 531320 604
rect 531372 592 531378 604
rect 532234 592 532240 604
rect 531372 564 532240 592
rect 531372 552 531378 564
rect 532234 552 532240 564
rect 532292 552 532298 604
rect 538214 552 538220 604
rect 538272 592 538278 604
rect 539318 592 539324 604
rect 538272 564 539324 592
rect 538272 552 538278 564
rect 539318 552 539324 564
rect 539376 552 539382 604
rect 542354 552 542360 604
rect 542412 592 542418 604
rect 542906 592 542912 604
rect 542412 564 542912 592
rect 542412 552 542418 564
rect 542906 552 542912 564
rect 542964 552 542970 604
<< via1 >>
rect 315948 700816 316000 700868
rect 397460 700816 397512 700868
rect 325608 700748 325660 700800
rect 413652 700748 413704 700800
rect 333888 700680 333940 700732
rect 429844 700680 429896 700732
rect 342168 700612 342220 700664
rect 462320 700612 462372 700664
rect 351828 700544 351880 700596
rect 478512 700544 478564 700596
rect 360108 700476 360160 700528
rect 494796 700476 494848 700528
rect 289728 700408 289780 700460
rect 332508 700408 332560 700460
rect 368388 700408 368440 700460
rect 527180 700408 527232 700460
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 273168 700340 273220 700392
rect 283840 700340 283892 700392
rect 299388 700340 299440 700392
rect 348792 700340 348844 700392
rect 376668 700340 376720 700392
rect 543464 700340 543516 700392
rect 281448 700272 281500 700324
rect 300124 700272 300176 700324
rect 307668 700272 307720 700324
rect 364984 700272 365036 700324
rect 386328 700272 386380 700324
rect 559656 700272 559708 700324
rect 170312 700204 170364 700256
rect 171048 700204 171100 700256
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 89168 699660 89220 699712
rect 89628 699660 89680 699712
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 264888 699660 264940 699712
rect 267648 699660 267700 699712
rect 8024 698232 8076 698284
rect 8208 698232 8260 698284
rect 137744 698232 137796 698284
rect 137928 698232 137980 698284
rect 393964 696940 394016 696992
rect 580172 696940 580224 696992
rect 154120 695512 154172 695564
rect 154212 695512 154264 695564
rect 8208 695444 8260 695496
rect 137928 695444 137980 695496
rect 219164 695444 219216 695496
rect 72700 694084 72752 694136
rect 154212 688576 154264 688628
rect 154396 688576 154448 688628
rect 8116 685899 8168 685908
rect 8116 685865 8125 685899
rect 8125 685865 8159 685899
rect 8159 685865 8168 685899
rect 8116 685856 8168 685865
rect 137836 685899 137888 685908
rect 137836 685865 137845 685899
rect 137845 685865 137879 685899
rect 137879 685865 137888 685899
rect 137836 685856 137888 685865
rect 219072 685899 219124 685908
rect 219072 685865 219081 685899
rect 219081 685865 219115 685899
rect 219115 685865 219124 685899
rect 219072 685856 219124 685865
rect 392584 685856 392636 685908
rect 580172 685856 580224 685908
rect 154396 685788 154448 685840
rect 72516 684607 72568 684616
rect 72516 684573 72525 684607
rect 72525 684573 72559 684607
rect 72559 684573 72568 684607
rect 72516 684564 72568 684573
rect 72516 684428 72568 684480
rect 3332 681708 3384 681760
rect 6184 681708 6236 681760
rect 8116 678988 8168 679040
rect 137836 678988 137888 679040
rect 8024 678920 8076 678972
rect 137744 678920 137796 678972
rect 154304 676243 154356 676252
rect 154304 676209 154313 676243
rect 154313 676209 154347 676243
rect 154347 676209 154356 676243
rect 154304 676200 154356 676209
rect 218980 676175 219032 676184
rect 218980 676141 218989 676175
rect 218989 676141 219023 676175
rect 219023 676141 219032 676175
rect 218980 676132 219032 676141
rect 72792 676107 72844 676116
rect 72792 676073 72801 676107
rect 72801 676073 72835 676107
rect 72835 676073 72844 676107
rect 72792 676064 72844 676073
rect 8024 673480 8076 673532
rect 8208 673480 8260 673532
rect 137744 673480 137796 673532
rect 137928 673480 137980 673532
rect 154304 673480 154356 673532
rect 154488 673480 154540 673532
rect 72792 669332 72844 669384
rect 72792 669196 72844 669248
rect 219072 666544 219124 666596
rect 72884 659608 72936 659660
rect 73068 659608 73120 659660
rect 219164 659608 219216 659660
rect 219348 659608 219400 659660
rect 73068 656820 73120 656872
rect 219348 656820 219400 656872
rect 8024 654100 8076 654152
rect 8208 654100 8260 654152
rect 137744 654100 137796 654152
rect 137928 654100 137980 654152
rect 154304 654100 154356 654152
rect 154488 654100 154540 654152
rect 72976 647275 73028 647284
rect 72976 647241 72985 647275
rect 72985 647241 73019 647275
rect 73019 647241 73028 647275
rect 72976 647232 73028 647241
rect 219256 647275 219308 647284
rect 219256 647241 219265 647275
rect 219265 647241 219299 647275
rect 219299 647241 219308 647275
rect 219256 647232 219308 647241
rect 72976 640364 73028 640416
rect 219256 640364 219308 640416
rect 72792 640228 72844 640280
rect 219072 640228 219124 640280
rect 398104 638936 398156 638988
rect 579896 638936 579948 638988
rect 72792 637508 72844 637560
rect 72884 637508 72936 637560
rect 219072 637508 219124 637560
rect 219164 637508 219216 637560
rect 8024 634788 8076 634840
rect 8208 634788 8260 634840
rect 137744 634788 137796 634840
rect 137928 634788 137980 634840
rect 154304 634788 154356 634840
rect 154488 634788 154540 634840
rect 73068 626535 73120 626544
rect 73068 626501 73077 626535
rect 73077 626501 73111 626535
rect 73111 626501 73120 626535
rect 73068 626492 73120 626501
rect 219348 626535 219400 626544
rect 219348 626501 219357 626535
rect 219357 626501 219391 626535
rect 219391 626501 219400 626535
rect 219348 626492 219400 626501
rect 3056 623772 3108 623824
rect 133144 623772 133196 623824
rect 73068 616879 73120 616888
rect 73068 616845 73077 616879
rect 73077 616845 73111 616879
rect 73111 616845 73120 616879
rect 73068 616836 73120 616845
rect 219348 616879 219400 616888
rect 219348 616845 219357 616879
rect 219357 616845 219391 616879
rect 219391 616845 219400 616879
rect 219348 616836 219400 616845
rect 8024 615476 8076 615528
rect 8208 615476 8260 615528
rect 137744 615476 137796 615528
rect 137928 615476 137980 615528
rect 154304 615476 154356 615528
rect 154488 615476 154540 615528
rect 73068 611396 73120 611448
rect 219348 611396 219400 611448
rect 72884 611260 72936 611312
rect 219072 608719 219124 608728
rect 219072 608685 219081 608719
rect 219081 608685 219115 608719
rect 219115 608685 219124 608719
rect 219072 608676 219124 608685
rect 219072 608540 219124 608592
rect 72976 601536 73028 601588
rect 73160 601536 73212 601588
rect 219256 601579 219308 601588
rect 219256 601545 219265 601579
rect 219265 601545 219299 601579
rect 219299 601545 219308 601579
rect 219256 601536 219308 601545
rect 72976 598884 73028 598936
rect 219256 598884 219308 598936
rect 8024 596164 8076 596216
rect 8208 596164 8260 596216
rect 137744 596164 137796 596216
rect 137928 596164 137980 596216
rect 154304 596164 154356 596216
rect 154488 596164 154540 596216
rect 392676 592016 392728 592068
rect 580172 592016 580224 592068
rect 72884 589339 72936 589348
rect 72884 589305 72893 589339
rect 72893 589305 72927 589339
rect 72927 589305 72936 589339
rect 72884 589296 72936 589305
rect 219164 589339 219216 589348
rect 219164 589305 219173 589339
rect 219173 589305 219207 589339
rect 219207 589305 219216 589339
rect 219164 589296 219216 589305
rect 8024 589271 8076 589280
rect 8024 589237 8033 589271
rect 8033 589237 8067 589271
rect 8067 589237 8076 589271
rect 8024 589228 8076 589237
rect 137744 589271 137796 589280
rect 137744 589237 137753 589271
rect 137753 589237 137787 589271
rect 137787 589237 137796 589271
rect 137744 589228 137796 589237
rect 154304 589271 154356 589280
rect 154304 589237 154313 589271
rect 154313 589237 154347 589271
rect 154347 589237 154356 589271
rect 154304 589228 154356 589237
rect 72700 582360 72752 582412
rect 72884 582360 72936 582412
rect 218980 582360 219032 582412
rect 219164 582360 219216 582412
rect 8024 579751 8076 579760
rect 8024 579717 8033 579751
rect 8033 579717 8067 579751
rect 8067 579717 8076 579751
rect 8024 579708 8076 579717
rect 137744 579751 137796 579760
rect 137744 579717 137753 579751
rect 137753 579717 137787 579751
rect 137787 579717 137796 579751
rect 137744 579708 137796 579717
rect 154304 579751 154356 579760
rect 154304 579717 154313 579751
rect 154313 579717 154347 579751
rect 154347 579717 154356 579751
rect 154304 579708 154356 579717
rect 7932 579572 7984 579624
rect 8116 579572 8168 579624
rect 72700 579572 72752 579624
rect 137652 579572 137704 579624
rect 154212 579572 154264 579624
rect 154396 579572 154448 579624
rect 218980 579572 219032 579624
rect 72608 569959 72660 569968
rect 72608 569925 72617 569959
rect 72617 569925 72651 569959
rect 72651 569925 72660 569959
rect 72608 569916 72660 569925
rect 137560 569959 137612 569968
rect 137560 569925 137569 569959
rect 137569 569925 137603 569959
rect 137603 569925 137612 569959
rect 137560 569916 137612 569925
rect 218888 569959 218940 569968
rect 218888 569925 218897 569959
rect 218897 569925 218931 569959
rect 218931 569925 218940 569959
rect 218888 569916 218940 569925
rect 4068 567196 4120 567248
rect 15844 567196 15896 567248
rect 72608 563048 72660 563100
rect 137560 563048 137612 563100
rect 218888 563048 218940 563100
rect 7932 562912 7984 562964
rect 8116 562912 8168 562964
rect 72700 562912 72752 562964
rect 137652 562912 137704 562964
rect 154212 562912 154264 562964
rect 154396 562912 154448 562964
rect 218980 562912 219032 562964
rect 137652 560235 137704 560244
rect 137652 560201 137661 560235
rect 137661 560201 137695 560235
rect 137695 560201 137704 560235
rect 137652 560192 137704 560201
rect 72608 553435 72660 553444
rect 72608 553401 72617 553435
rect 72617 553401 72651 553435
rect 72651 553401 72660 553435
rect 72608 553392 72660 553401
rect 218888 553435 218940 553444
rect 218888 553401 218897 553435
rect 218897 553401 218931 553435
rect 218931 553401 218940 553435
rect 218888 553392 218940 553401
rect 72608 550647 72660 550656
rect 72608 550613 72617 550647
rect 72617 550613 72651 550647
rect 72651 550613 72660 550647
rect 72608 550604 72660 550613
rect 137836 550604 137888 550656
rect 218888 550647 218940 550656
rect 218888 550613 218897 550647
rect 218897 550613 218931 550647
rect 218931 550613 218940 550647
rect 218888 550604 218940 550613
rect 8024 550579 8076 550588
rect 8024 550545 8033 550579
rect 8033 550545 8067 550579
rect 8067 550545 8076 550579
rect 8024 550536 8076 550545
rect 396724 545096 396776 545148
rect 580172 545096 580224 545148
rect 72608 543736 72660 543788
rect 218888 543736 218940 543788
rect 72700 543600 72752 543652
rect 137652 543600 137704 543652
rect 137836 543600 137888 543652
rect 218980 543600 219032 543652
rect 8208 540948 8260 541000
rect 72608 534123 72660 534132
rect 72608 534089 72617 534123
rect 72617 534089 72651 534123
rect 72651 534089 72660 534123
rect 72608 534080 72660 534089
rect 137652 534012 137704 534064
rect 137836 534012 137888 534064
rect 72608 531335 72660 531344
rect 72608 531301 72617 531335
rect 72617 531301 72651 531335
rect 72651 531301 72660 531335
rect 72608 531292 72660 531301
rect 154396 531267 154448 531276
rect 154396 531233 154405 531267
rect 154405 531233 154439 531267
rect 154439 531233 154448 531267
rect 154396 531224 154448 531233
rect 72700 524288 72752 524340
rect 72884 524288 72936 524340
rect 218980 524288 219032 524340
rect 219164 524288 219216 524340
rect 8208 521636 8260 521688
rect 8392 521636 8444 521688
rect 137928 521636 137980 521688
rect 138112 521636 138164 521688
rect 154488 521636 154540 521688
rect 154396 511955 154448 511964
rect 154396 511921 154405 511955
rect 154405 511921 154439 511955
rect 154439 511921 154448 511955
rect 154396 511912 154448 511921
rect 3332 509736 3384 509788
rect 10324 509736 10376 509788
rect 8208 502324 8260 502376
rect 8392 502324 8444 502376
rect 72608 502324 72660 502376
rect 73068 502324 73120 502376
rect 137928 502324 137980 502376
rect 138112 502324 138164 502376
rect 154488 502324 154540 502376
rect 218888 502324 218940 502376
rect 219348 502324 219400 502376
rect 392768 498176 392820 498228
rect 579988 498176 580040 498228
rect 137652 492600 137704 492652
rect 137836 492600 137888 492652
rect 154212 492600 154264 492652
rect 154396 492600 154448 492652
rect 8116 485800 8168 485852
rect 400864 485800 400916 485852
rect 579988 485800 580040 485852
rect 8208 485732 8260 485784
rect 7932 482944 7984 482996
rect 8208 482944 8260 482996
rect 72884 480224 72936 480276
rect 73068 480224 73120 480276
rect 219164 480224 219216 480276
rect 219348 480224 219400 480276
rect 8116 466420 8168 466472
rect 137744 466488 137796 466540
rect 154304 466420 154356 466472
rect 154488 466420 154540 466472
rect 8208 466352 8260 466404
rect 137652 466352 137704 466404
rect 137376 463632 137428 463684
rect 137652 463632 137704 463684
rect 395344 462340 395396 462392
rect 579988 462340 580040 462392
rect 72884 460912 72936 460964
rect 73068 460912 73120 460964
rect 219164 460912 219216 460964
rect 219348 460912 219400 460964
rect 8024 453976 8076 454028
rect 154304 453976 154356 454028
rect 3332 451392 3384 451444
rect 11704 451392 11756 451444
rect 399484 451256 399536 451308
rect 579988 451256 580040 451308
rect 137560 447108 137612 447160
rect 137652 447040 137704 447092
rect 7932 444431 7984 444440
rect 7932 444397 7941 444431
rect 7941 444397 7975 444431
rect 7975 444397 7984 444431
rect 7932 444388 7984 444397
rect 154212 444431 154264 444440
rect 154212 444397 154221 444431
rect 154221 444397 154255 444431
rect 154255 444397 154264 444431
rect 154212 444388 154264 444397
rect 72976 444320 73028 444372
rect 73160 444320 73212 444372
rect 219256 444320 219308 444372
rect 219440 444320 219492 444372
rect 3332 437656 3384 437708
rect 4804 437656 4856 437708
rect 8024 427796 8076 427848
rect 137744 427796 137796 427848
rect 154304 427796 154356 427848
rect 8116 427728 8168 427780
rect 137836 427728 137888 427780
rect 154396 427728 154448 427780
rect 7840 425008 7892 425060
rect 8116 425008 8168 425060
rect 137560 425008 137612 425060
rect 137836 425008 137888 425060
rect 154120 425008 154172 425060
rect 154396 425008 154448 425060
rect 72700 418208 72752 418260
rect 218980 418208 219032 418260
rect 72608 418072 72660 418124
rect 218888 418072 218940 418124
rect 392860 415420 392912 415472
rect 580080 415420 580132 415472
rect 263600 415352 263652 415404
rect 264888 415352 264940 415404
rect 298376 415352 298428 415404
rect 299388 415352 299440 415404
rect 359280 415352 359332 415404
rect 360108 415352 360160 415404
rect 385316 415352 385368 415404
rect 386328 415352 386380 415404
rect 154304 415148 154356 415200
rect 220176 415148 220228 415200
rect 137744 415080 137796 415132
rect 211436 415080 211488 415132
rect 350540 415080 350592 415132
rect 351828 415080 351880 415132
rect 106188 415012 106240 415064
rect 202420 415012 202472 415064
rect 89628 414944 89680 414996
rect 194048 414944 194100 414996
rect 72608 414876 72660 414928
rect 185400 414876 185452 414928
rect 41328 414808 41380 414860
rect 176660 414808 176712 414860
rect 218888 414808 218940 414860
rect 246212 414808 246264 414860
rect 24768 414740 24820 414792
rect 168012 414740 168064 414792
rect 202788 414740 202840 414792
rect 237564 414740 237616 414792
rect 8024 414672 8076 414724
rect 159364 414672 159416 414724
rect 171048 414672 171100 414724
rect 228824 414672 228876 414724
rect 235908 414672 235960 414724
rect 254952 414672 255004 414724
rect 272340 414672 272392 414724
rect 273168 414672 273220 414724
rect 324504 414196 324556 414248
rect 325608 414196 325660 414248
rect 579896 412564 579948 412616
rect 580264 412564 580316 412616
rect 3516 409776 3568 409828
rect 151820 409776 151872 409828
rect 391940 409232 391992 409284
rect 393964 409232 394016 409284
rect 393964 404336 394016 404388
rect 580080 404336 580132 404388
rect 3424 404268 3476 404320
rect 152372 404268 152424 404320
rect 6184 398760 6236 398812
rect 153108 398760 153160 398812
rect 391940 398760 391992 398812
rect 580080 398760 580132 398812
rect 391940 394612 391992 394664
rect 580356 394612 580408 394664
rect 3700 393252 3752 393304
rect 153108 393252 153160 393304
rect 391940 389104 391992 389156
rect 398104 389104 398156 389156
rect 3608 386316 3660 386368
rect 153108 386316 153160 386368
rect 391940 383596 391992 383648
rect 580448 383596 580500 383648
rect 133144 380808 133196 380860
rect 152556 380808 152608 380860
rect 391940 378088 391992 378140
rect 580540 378088 580592 378140
rect 3884 375300 3936 375352
rect 152556 375300 152608 375352
rect 3792 369792 3844 369844
rect 152924 369792 152976 369844
rect 392584 368500 392636 368552
rect 580080 368500 580132 368552
rect 391940 367004 391992 367056
rect 580632 367004 580684 367056
rect 15844 364284 15896 364336
rect 153108 364284 153160 364336
rect 391940 362856 391992 362908
rect 580724 362856 580776 362908
rect 4068 358708 4120 358760
rect 153108 358708 153160 358760
rect 392676 357416 392728 357468
rect 580080 357416 580132 357468
rect 391940 357348 391992 357400
rect 396724 357348 396776 357400
rect 3976 353200 4028 353252
rect 153108 353200 153160 353252
rect 391940 351840 391992 351892
rect 580816 351840 580868 351892
rect 10324 347692 10376 347744
rect 152924 347692 152976 347744
rect 391940 346332 391992 346384
rect 580908 346332 580960 346384
rect 3332 342184 3384 342236
rect 152556 342184 152608 342236
rect 4804 336676 4856 336728
rect 153108 336676 153160 336728
rect 391940 336676 391992 336728
rect 400864 336676 400916 336728
rect 11704 331168 11756 331220
rect 153108 331168 153160 331220
rect 391940 330352 391992 330404
rect 395344 330352 395396 330404
rect 391940 325592 391992 325644
rect 399484 325592 399536 325644
rect 3608 324232 3660 324284
rect 153108 324232 153160 324284
rect 579896 322736 579948 322788
rect 580172 322736 580224 322788
rect 392768 321580 392820 321632
rect 580172 321580 580224 321632
rect 391940 320084 391992 320136
rect 579896 320084 579948 320136
rect 3516 318724 3568 318776
rect 153108 318724 153160 318776
rect 3424 313216 3476 313268
rect 152372 313216 152424 313268
rect 392860 310496 392912 310548
rect 579620 310496 579672 310548
rect 391940 309544 391992 309596
rect 393964 309544 394016 309596
rect 3056 307708 3108 307760
rect 152556 307708 152608 307760
rect 391940 304920 391992 304972
rect 580264 304920 580316 304972
rect 3792 302132 3844 302184
rect 153108 302132 153160 302184
rect 3700 296624 3752 296676
rect 152740 296624 152792 296676
rect 3424 289824 3476 289876
rect 152188 289824 152240 289876
rect 391940 288328 391992 288380
rect 580356 288328 580408 288380
rect 2964 284316 3016 284368
rect 152004 284316 152056 284368
rect 3516 280100 3568 280152
rect 152924 280100 152976 280152
rect 392584 274660 392636 274712
rect 580172 274660 580224 274712
rect 391940 273164 391992 273216
rect 580264 273164 580316 273216
rect 3516 267724 3568 267776
rect 153108 267724 153160 267776
rect 391940 263576 391992 263628
rect 579804 263576 579856 263628
rect 3424 262216 3476 262268
rect 153108 262216 153160 262268
rect 391940 252492 391992 252544
rect 579804 252492 579856 252544
rect 3424 249772 3476 249824
rect 153108 249772 153160 249824
rect 3700 233248 3752 233300
rect 153108 233248 153160 233300
rect 392768 229032 392820 229084
rect 580172 229032 580224 229084
rect 3516 223524 3568 223576
rect 152464 223524 152516 223576
rect 392676 217948 392728 218000
rect 580172 217948 580224 218000
rect 3608 216656 3660 216708
rect 153016 216656 153068 216708
rect 391940 208360 391992 208412
rect 395344 208360 395396 208412
rect 3148 208292 3200 208344
rect 152556 208292 152608 208344
rect 392584 205572 392636 205624
rect 579804 205572 579856 205624
rect 3516 200132 3568 200184
rect 152004 200132 152056 200184
rect 3424 182180 3476 182232
rect 152464 182180 152516 182232
rect 392492 182112 392544 182164
rect 580172 182112 580224 182164
rect 3056 180752 3108 180804
rect 152648 180752 152700 180804
rect 391940 176672 391992 176724
rect 519084 176672 519136 176724
rect 188068 173995 188120 174004
rect 188068 173961 188077 173995
rect 188077 173961 188111 173995
rect 188111 173961 188120 173995
rect 188068 173952 188120 173961
rect 211068 173816 211120 173868
rect 219348 173748 219400 173800
rect 243268 173816 243320 173868
rect 246304 173816 246356 173868
rect 253848 173816 253900 173868
rect 320456 173816 320508 173868
rect 409880 173816 409932 173868
rect 241888 173748 241940 173800
rect 246948 173748 247000 173800
rect 254308 173748 254360 173800
rect 323308 173748 323360 173800
rect 416780 173748 416832 173800
rect 122748 173680 122800 173732
rect 204076 173680 204128 173732
rect 213828 173680 213880 173732
rect 240876 173680 240928 173732
rect 245568 173680 245620 173732
rect 253388 173680 253440 173732
rect 326160 173680 326212 173732
rect 425060 173680 425112 173732
rect 118608 173612 118660 173664
rect 202604 173612 202656 173664
rect 239956 173612 240008 173664
rect 242808 173612 242860 173664
rect 252376 173612 252428 173664
rect 329012 173612 329064 173664
rect 431960 173612 432012 173664
rect 111708 173544 111760 173596
rect 199752 173544 199804 173596
rect 206928 173544 206980 173596
rect 235172 173544 235224 173596
rect 244924 173544 244976 173596
rect 252928 173544 252980 173596
rect 331956 173544 332008 173596
rect 438860 173544 438912 173596
rect 35164 173476 35216 173528
rect 168104 173476 168156 173528
rect 204168 173476 204220 173528
rect 241428 173476 241480 173528
rect 251916 173476 251968 173528
rect 334808 173476 334860 173528
rect 445760 173476 445812 173528
rect 29644 173408 29696 173460
rect 165252 173408 165304 173460
rect 201408 173408 201460 173460
rect 19984 173340 20036 173392
rect 161388 173340 161440 173392
rect 202788 173340 202840 173392
rect 235264 173408 235316 173460
rect 248052 173408 248104 173460
rect 248328 173408 248380 173460
rect 254768 173408 254820 173460
rect 337660 173408 337712 173460
rect 452660 173408 452712 173460
rect 235632 173340 235684 173392
rect 238668 173340 238720 173392
rect 250996 173340 251048 173392
rect 312544 173340 312596 173392
rect 28264 173272 28316 173324
rect 164792 173272 164844 173324
rect 200028 173272 200080 173324
rect 235908 173272 235960 173324
rect 249524 173272 249576 173324
rect 273444 173272 273496 173324
rect 287704 173272 287756 173324
rect 18604 173204 18656 173256
rect 160928 173204 160980 173256
rect 197268 173204 197320 173256
rect 237104 173204 237156 173256
rect 237288 173204 237340 173256
rect 250536 173204 250588 173256
rect 262496 173204 262548 173256
rect 266544 173204 266596 173256
rect 281172 173204 281224 173256
rect 288348 173204 288400 173256
rect 10324 173136 10376 173188
rect 157616 173136 157668 173188
rect 194416 173136 194468 173188
rect 232780 173136 232832 173188
rect 249064 173136 249116 173188
rect 251088 173136 251140 173188
rect 255780 173136 255832 173188
rect 263876 173136 263928 173188
rect 267004 173136 267056 173188
rect 317512 173204 317564 173256
rect 217876 173068 217928 173120
rect 242348 173068 242400 173120
rect 261944 173068 261996 173120
rect 265256 173068 265308 173120
rect 267740 173068 267792 173120
rect 268936 173068 268988 173120
rect 274916 173068 274968 173120
rect 275836 173068 275888 173120
rect 277768 173068 277820 173120
rect 278688 173068 278740 173120
rect 280712 173068 280764 173120
rect 281356 173068 281408 173120
rect 281632 173068 281684 173120
rect 282828 173068 282880 173120
rect 340512 173340 340564 173392
rect 459560 173340 459612 173392
rect 324688 173204 324740 173256
rect 325608 173204 325660 173256
rect 325700 173204 325752 173256
rect 326896 173204 326948 173256
rect 331312 173272 331364 173324
rect 343456 173272 343508 173324
rect 467840 173272 467892 173324
rect 330484 173204 330536 173256
rect 331128 173204 331180 173256
rect 333336 173204 333388 173256
rect 333888 173204 333940 173256
rect 337200 173204 337252 173256
rect 337936 173204 337988 173256
rect 338580 173204 338632 173256
rect 339224 173204 339276 173256
rect 340052 173204 340104 173256
rect 340696 173204 340748 173256
rect 349160 173204 349212 173256
rect 327632 173136 327684 173188
rect 328368 173136 328420 173188
rect 328552 173136 328604 173188
rect 329656 173136 329708 173188
rect 330024 173136 330076 173188
rect 330944 173136 330996 173188
rect 331404 173136 331456 173188
rect 332416 173136 332468 173188
rect 332876 173136 332928 173188
rect 333704 173136 333756 173188
rect 335728 173136 335780 173188
rect 336556 173136 336608 173188
rect 336740 173136 336792 173188
rect 338028 173136 338080 173188
rect 338120 173136 338172 173188
rect 339316 173136 339368 173188
rect 339592 173136 339644 173188
rect 340788 173136 340840 173188
rect 342444 173136 342496 173188
rect 343548 173136 343600 173188
rect 343916 173136 343968 173188
rect 344836 173136 344888 173188
rect 345296 173136 345348 173188
rect 346308 173136 346360 173188
rect 346768 173136 346820 173188
rect 347596 173136 347648 173188
rect 348240 173136 348292 173188
rect 349068 173136 349120 173188
rect 350632 173136 350684 173188
rect 351736 173136 351788 173188
rect 352012 173136 352064 173188
rect 353208 173136 353260 173188
rect 474740 173204 474792 173256
rect 481640 173136 481692 173188
rect 519084 173136 519136 173188
rect 580264 173136 580316 173188
rect 402980 173068 403032 173120
rect 214564 173000 214616 173052
rect 216496 173000 216548 173052
rect 216588 173000 216640 173052
rect 244740 173000 244792 173052
rect 249708 173000 249760 173052
rect 255320 173000 255372 173052
rect 314660 173000 314712 173052
rect 396080 173000 396132 173052
rect 227628 172932 227680 172984
rect 246212 172932 246264 172984
rect 270592 172932 270644 172984
rect 271604 172932 271656 172984
rect 272064 172932 272116 172984
rect 272984 172932 273036 172984
rect 310336 172932 310388 172984
rect 385408 172932 385460 172984
rect 223488 172864 223540 172916
rect 234252 172864 234304 172916
rect 234528 172864 234580 172916
rect 247592 172864 247644 172916
rect 279240 172864 279292 172916
rect 279976 172864 280028 172916
rect 307484 172864 307536 172916
rect 229008 172796 229060 172848
rect 246672 172796 246724 172848
rect 346400 172796 346452 172848
rect 354864 172796 354916 172848
rect 355968 172796 356020 172848
rect 356336 172796 356388 172848
rect 357348 172796 357400 172848
rect 357808 172796 357860 172848
rect 358728 172796 358780 172848
rect 359188 172796 359240 172848
rect 360108 172796 360160 172848
rect 360660 172796 360712 172848
rect 361488 172796 361540 172848
rect 361580 172796 361632 172848
rect 362776 172796 362828 172848
rect 363052 172796 363104 172848
rect 364064 172796 364116 172848
rect 364524 172796 364576 172848
rect 365444 172796 365496 172848
rect 365904 172796 365956 172848
rect 366916 172796 366968 172848
rect 367376 172796 367428 172848
rect 368296 172796 368348 172848
rect 368756 172796 368808 172848
rect 369676 172796 369728 172848
rect 370228 172796 370280 172848
rect 371056 172796 371108 172848
rect 371700 172796 371752 172848
rect 372528 172796 372580 172848
rect 372620 172796 372672 172848
rect 373908 172796 373960 172848
rect 232504 172728 232556 172780
rect 245200 172728 245252 172780
rect 256608 172728 256660 172780
rect 258172 172728 258224 172780
rect 265348 172728 265400 172780
rect 266176 172728 266228 172780
rect 266820 172728 266872 172780
rect 267648 172728 267700 172780
rect 268200 172728 268252 172780
rect 269028 172728 269080 172780
rect 269212 172728 269264 172780
rect 270224 172728 270276 172780
rect 276388 172728 276440 172780
rect 277124 172728 277176 172780
rect 321836 172728 321888 172780
rect 322848 172728 322900 172780
rect 340972 172728 341024 172780
rect 342076 172728 342128 172780
rect 353484 172728 353536 172780
rect 354496 172728 354548 172780
rect 354772 172728 354824 172780
rect 355416 172728 355468 172780
rect 360200 172728 360252 172780
rect 361396 172728 361448 172780
rect 373080 172728 373132 172780
rect 373816 172728 373868 172780
rect 374092 172864 374144 172916
rect 375196 172864 375248 172916
rect 375472 172864 375524 172916
rect 376576 172864 376628 172916
rect 376944 172864 376996 172916
rect 377956 172864 378008 172916
rect 378416 172864 378468 172916
rect 379336 172864 379388 172916
rect 374552 172796 374604 172848
rect 375104 172796 375156 172848
rect 378324 172728 378376 172780
rect 231124 172660 231176 172712
rect 243084 172660 243136 172712
rect 243544 172660 243596 172712
rect 253848 172660 253900 172712
rect 256700 172660 256752 172712
rect 236644 172592 236696 172644
rect 255228 172592 255280 172644
rect 257712 172592 257764 172644
rect 261484 172592 261536 172644
rect 262864 172592 262916 172644
rect 262956 172592 263008 172644
rect 264244 172592 264296 172644
rect 265808 172592 265860 172644
rect 268384 172592 268436 172644
rect 275376 172592 275428 172644
rect 278044 172592 278096 172644
rect 278780 172592 278832 172644
rect 280068 172592 280120 172644
rect 280160 172592 280212 172644
rect 281448 172592 281500 172644
rect 283564 172592 283616 172644
rect 290464 172592 290516 172644
rect 291200 172592 291252 172644
rect 292396 172592 292448 172644
rect 292672 172592 292724 172644
rect 293776 172592 293828 172644
rect 294512 172592 294564 172644
rect 295248 172592 295300 172644
rect 295524 172592 295576 172644
rect 296536 172592 296588 172644
rect 296996 172592 297048 172644
rect 297916 172592 297968 172644
rect 298836 172592 298888 172644
rect 299388 172592 299440 172644
rect 299848 172592 299900 172644
rect 300584 172592 300636 172644
rect 302700 172592 302752 172644
rect 303344 172592 303396 172644
rect 305552 172592 305604 172644
rect 306104 172592 306156 172644
rect 307024 172592 307076 172644
rect 307576 172592 307628 172644
rect 327080 172592 327132 172644
rect 328184 172592 328236 172644
rect 334348 172592 334400 172644
rect 335176 172592 335228 172644
rect 383660 172592 383712 172644
rect 384948 172592 385000 172644
rect 385040 172592 385092 172644
rect 386328 172592 386380 172644
rect 386512 172592 386564 172644
rect 387708 172592 387760 172644
rect 387984 172592 388036 172644
rect 389088 172592 389140 172644
rect 389364 172592 389416 172644
rect 390468 172592 390520 172644
rect 215944 172524 215996 172576
rect 217968 172524 218020 172576
rect 238024 172524 238076 172576
rect 243544 172524 243596 172576
rect 248604 172524 248656 172576
rect 254584 172524 254636 172576
rect 256240 172524 256292 172576
rect 260104 172524 260156 172576
rect 260932 172524 260984 172576
rect 261024 172524 261076 172576
rect 262128 172524 262180 172576
rect 283104 172524 283156 172576
rect 284208 172524 284260 172576
rect 284484 172524 284536 172576
rect 285496 172524 285548 172576
rect 285956 172524 286008 172576
rect 286968 172524 287020 172576
rect 287336 172524 287388 172576
rect 288348 172524 288400 172576
rect 288808 172524 288860 172576
rect 289728 172524 289780 172576
rect 290280 172524 290332 172576
rect 291108 172524 291160 172576
rect 291660 172524 291712 172576
rect 292488 172524 292540 172576
rect 293132 172524 293184 172576
rect 293868 172524 293920 172576
rect 294052 172524 294104 172576
rect 295064 172524 295116 172576
rect 295984 172524 296036 172576
rect 296628 172524 296680 172576
rect 297456 172524 297508 172576
rect 298008 172524 298060 172576
rect 298376 172524 298428 172576
rect 299204 172524 299256 172576
rect 300308 172524 300360 172576
rect 300768 172524 300820 172576
rect 301228 172524 301280 172576
rect 302056 172524 302108 172576
rect 302240 172524 302292 172576
rect 303436 172524 303488 172576
rect 303620 172524 303672 172576
rect 304816 172524 304868 172576
rect 305092 172524 305144 172576
rect 306196 172524 306248 172576
rect 306564 172524 306616 172576
rect 307668 172524 307720 172576
rect 307944 172524 307996 172576
rect 308956 172524 309008 172576
rect 309416 172524 309468 172576
rect 310428 172524 310480 172576
rect 310796 172524 310848 172576
rect 311716 172524 311768 172576
rect 313280 172524 313332 172576
rect 314568 172524 314620 172576
rect 315120 172524 315172 172576
rect 315856 172524 315908 172576
rect 316132 172524 316184 172576
rect 317328 172524 317380 172576
rect 318984 172524 319036 172576
rect 320088 172524 320140 172576
rect 379796 172524 379848 172576
rect 380716 172524 380768 172576
rect 381268 172524 381320 172576
rect 382096 172524 382148 172576
rect 382648 172524 382700 172576
rect 383568 172524 383620 172576
rect 384120 172524 384172 172576
rect 384856 172524 384908 172576
rect 385592 172524 385644 172576
rect 386236 172524 386288 172576
rect 386972 172524 387024 172576
rect 387616 172524 387668 172576
rect 388444 172524 388496 172576
rect 388996 172524 389048 172576
rect 163504 172499 163556 172508
rect 163504 172465 163513 172499
rect 163513 172465 163547 172499
rect 163547 172465 163556 172499
rect 163504 172456 163556 172465
rect 185124 172456 185176 172508
rect 185400 172456 185452 172508
rect 224224 172456 224276 172508
rect 126888 171844 126940 171896
rect 205916 171844 205968 171896
rect 114468 171776 114520 171828
rect 200672 171776 200724 171828
rect 349620 171776 349672 171828
rect 483020 171776 483072 171828
rect 225512 171096 225564 171148
rect 226064 171096 226116 171148
rect 154580 171028 154632 171080
rect 155316 171028 155368 171080
rect 169760 171028 169812 171080
rect 170588 171028 170640 171080
rect 171140 171028 171192 171080
rect 172060 171028 172112 171080
rect 175372 171028 175424 171080
rect 175924 171028 175976 171080
rect 176660 171028 176712 171080
rect 177120 171028 177172 171080
rect 178040 171028 178092 171080
rect 178316 171028 178368 171080
rect 179420 171028 179472 171080
rect 179880 171028 179932 171080
rect 186412 171028 186464 171080
rect 186964 171028 187016 171080
rect 187792 171028 187844 171080
rect 188436 171028 188488 171080
rect 189080 171028 189132 171080
rect 189356 171028 189408 171080
rect 190552 171028 190604 171080
rect 191196 171028 191248 171080
rect 191932 171028 191984 171080
rect 192668 171028 192720 171080
rect 193312 171028 193364 171080
rect 194140 171028 194192 171080
rect 194692 171028 194744 171080
rect 195612 171028 195664 171080
rect 202972 171028 203024 171080
rect 203156 171028 203208 171080
rect 204260 171028 204312 171080
rect 205180 171028 205232 171080
rect 208400 171028 208452 171080
rect 209044 171028 209096 171080
rect 211252 171028 211304 171080
rect 211804 171028 211856 171080
rect 214012 171028 214064 171080
rect 214748 171028 214800 171080
rect 227812 171028 227864 171080
rect 228548 171028 228600 171080
rect 229192 171028 229244 171080
rect 230020 171028 230072 171080
rect 230480 171028 230532 171080
rect 230940 171028 230992 171080
rect 237472 171028 237524 171080
rect 238116 171028 238168 171080
rect 240508 171028 240560 171080
rect 241152 171028 241204 171080
rect 393228 171028 393280 171080
rect 579896 171028 579948 171080
rect 175280 170960 175332 171012
rect 175556 170960 175608 171012
rect 176752 170960 176804 171012
rect 177396 170960 177448 171012
rect 179512 170960 179564 171012
rect 180156 170960 180208 171012
rect 186320 170960 186372 171012
rect 186596 170960 186648 171012
rect 189172 170960 189224 171012
rect 189908 170960 189960 171012
rect 230572 170960 230624 171012
rect 231492 170960 231544 171012
rect 218060 170484 218112 170536
rect 218612 170484 218664 170536
rect 131028 170416 131080 170468
rect 207020 170416 207072 170468
rect 36544 170348 36596 170400
rect 169024 170348 169076 170400
rect 312268 170348 312320 170400
rect 390560 170348 390612 170400
rect 187700 169396 187752 169448
rect 188160 169396 188212 169448
rect 188160 169260 188212 169312
rect 159088 169124 159140 169176
rect 159272 169124 159324 169176
rect 137928 169056 137980 169108
rect 210240 169056 210292 169108
rect 217048 169056 217100 169108
rect 217232 169056 217284 169108
rect 96528 168988 96580 169040
rect 193496 168988 193548 169040
rect 350632 168988 350684 169040
rect 485780 168988 485832 169040
rect 157432 168308 157484 168360
rect 158260 168308 158312 168360
rect 158812 168308 158864 168360
rect 159732 168308 159784 168360
rect 212632 167900 212684 167952
rect 213276 167900 213328 167952
rect 194600 167832 194652 167884
rect 195060 167832 195112 167884
rect 142068 167696 142120 167748
rect 211712 167696 211764 167748
rect 32404 167628 32456 167680
rect 167644 167628 167696 167680
rect 178132 167628 178184 167680
rect 178868 167628 178920 167680
rect 352012 167628 352064 167680
rect 489920 167628 489972 167680
rect 209872 167424 209924 167476
rect 210332 167424 210384 167476
rect 207204 167356 207256 167408
rect 208032 167356 208084 167408
rect 156236 167016 156288 167068
rect 156880 167016 156932 167068
rect 201500 167016 201552 167068
rect 201684 167016 201736 167068
rect 215300 167016 215352 167068
rect 215484 167016 215536 167068
rect 256884 166948 256936 167000
rect 257068 166948 257120 167000
rect 133788 166336 133840 166388
rect 208492 166336 208544 166388
rect 38568 166268 38620 166320
rect 169944 166268 169996 166320
rect 353392 166268 353444 166320
rect 494060 166268 494112 166320
rect 3240 165520 3292 165572
rect 153108 165520 153160 165572
rect 174084 165316 174136 165368
rect 174544 165316 174596 165368
rect 144828 164840 144880 164892
rect 212724 164840 212776 164892
rect 354772 164840 354824 164892
rect 496820 164840 496872 164892
rect 181168 164228 181220 164280
rect 181720 164228 181772 164280
rect 182456 164228 182508 164280
rect 183192 164228 183244 164280
rect 183928 164228 183980 164280
rect 184480 164228 184532 164280
rect 168380 164160 168432 164212
rect 168656 164160 168708 164212
rect 172428 164160 172480 164212
rect 172704 164160 172756 164212
rect 206008 164203 206060 164212
rect 206008 164169 206017 164203
rect 206017 164169 206051 164203
rect 206051 164169 206060 164203
rect 206008 164160 206060 164169
rect 216956 164160 217008 164212
rect 217048 164160 217100 164212
rect 240508 164203 240560 164212
rect 240508 164169 240517 164203
rect 240517 164169 240551 164203
rect 240551 164169 240560 164203
rect 240508 164160 240560 164169
rect 256792 164160 256844 164212
rect 257068 164160 257120 164212
rect 385224 164203 385276 164212
rect 385224 164169 385233 164203
rect 385233 164169 385267 164203
rect 385267 164169 385276 164203
rect 385224 164160 385276 164169
rect 148968 163548 149020 163600
rect 214104 163548 214156 163600
rect 31024 163480 31076 163532
rect 165804 163480 165856 163532
rect 357164 163480 357216 163532
rect 500960 163480 501012 163532
rect 163044 162868 163096 162920
rect 223856 162911 223908 162920
rect 223856 162877 223865 162911
rect 223865 162877 223899 162911
rect 223899 162877 223908 162911
rect 223856 162868 223908 162877
rect 163136 162800 163188 162852
rect 163320 162800 163372 162852
rect 174084 162800 174136 162852
rect 174268 162800 174320 162852
rect 181168 162843 181220 162852
rect 181168 162809 181177 162843
rect 181177 162809 181211 162843
rect 181211 162809 181220 162843
rect 181168 162800 181220 162809
rect 151728 162188 151780 162240
rect 215392 162188 215444 162240
rect 21364 162120 21416 162172
rect 161572 162120 161624 162172
rect 201684 162120 201736 162172
rect 358544 162120 358596 162172
rect 503720 162120 503772 162172
rect 201684 161916 201736 161968
rect 163320 161372 163372 161424
rect 225420 161372 225472 161424
rect 132408 160760 132460 160812
rect 207112 160760 207164 160812
rect 55128 160692 55180 160744
rect 176844 160692 176896 160744
rect 360016 160692 360068 160744
rect 507860 160692 507912 160744
rect 201500 159400 201552 159452
rect 201868 159400 201920 159452
rect 128268 159332 128320 159384
rect 205732 159332 205784 159384
rect 361304 159332 361356 159384
rect 512000 159332 512052 159384
rect 393136 158652 393188 158704
rect 580172 158652 580224 158704
rect 146208 158040 146260 158092
rect 212632 158040 212684 158092
rect 11704 157972 11756 158024
rect 158904 157972 158956 158024
rect 198924 157496 198976 157548
rect 226524 157360 226576 157412
rect 226708 157360 226760 157412
rect 198924 157292 198976 157344
rect 385224 157335 385276 157344
rect 385224 157301 385233 157335
rect 385233 157301 385267 157335
rect 385267 157301 385276 157335
rect 385224 157292 385276 157301
rect 139308 156680 139360 156732
rect 209872 156680 209924 156732
rect 314384 156680 314436 156732
rect 393320 156680 393372 156732
rect 50988 156612 51040 156664
rect 175464 156612 175516 156664
rect 364064 156612 364116 156664
rect 516140 156612 516192 156664
rect 240508 156315 240560 156324
rect 240508 156281 240517 156315
rect 240517 156281 240551 156315
rect 240551 156281 240560 156315
rect 240508 156272 240560 156281
rect 150348 155252 150400 155304
rect 214012 155252 214064 155304
rect 315856 155252 315908 155304
rect 397460 155252 397512 155304
rect 42708 155184 42760 155236
rect 171416 155184 171468 155236
rect 365444 155184 365496 155236
rect 520280 155184 520332 155236
rect 206008 154615 206060 154624
rect 206008 154581 206017 154615
rect 206017 154581 206051 154615
rect 206051 154581 206060 154615
rect 206008 154572 206060 154581
rect 210056 154572 210108 154624
rect 210148 154572 210200 154624
rect 207204 154504 207256 154556
rect 207480 154504 207532 154556
rect 218244 154504 218296 154556
rect 218428 154504 218480 154556
rect 219532 154504 219584 154556
rect 219716 154504 219768 154556
rect 256976 154504 257028 154556
rect 257160 154504 257212 154556
rect 317144 153892 317196 153944
rect 400312 153892 400364 153944
rect 82728 153824 82780 153876
rect 188252 153824 188304 153876
rect 362684 153824 362736 153876
rect 513380 153824 513432 153876
rect 183928 153348 183980 153400
rect 183928 153212 183980 153264
rect 185216 153212 185268 153264
rect 185308 153212 185360 153264
rect 318616 152532 318668 152584
rect 404360 152532 404412 152584
rect 85488 152464 85540 152516
rect 189264 152464 189316 152516
rect 366824 152464 366876 152516
rect 524420 152464 524472 152516
rect 163044 151827 163096 151836
rect 163044 151793 163053 151827
rect 163053 151793 163087 151827
rect 163087 151793 163096 151827
rect 163044 151784 163096 151793
rect 225328 151827 225380 151836
rect 225328 151793 225337 151827
rect 225337 151793 225371 151827
rect 225371 151793 225380 151827
rect 225328 151784 225380 151793
rect 378140 151784 378192 151836
rect 378324 151784 378376 151836
rect 223764 151759 223816 151768
rect 223764 151725 223773 151759
rect 223773 151725 223807 151759
rect 223807 151725 223816 151759
rect 223764 151716 223816 151725
rect 319904 151104 319956 151156
rect 408500 151104 408552 151156
rect 89628 151036 89680 151088
rect 190644 151036 190696 151088
rect 279884 151036 279936 151088
rect 309140 151036 309192 151088
rect 368204 151036 368256 151088
rect 528560 151036 528612 151088
rect 321376 149744 321428 149796
rect 411260 149744 411312 149796
rect 92388 149676 92440 149728
rect 192024 149676 192076 149728
rect 369584 149676 369636 149728
rect 531320 149676 531372 149728
rect 322664 148384 322716 148436
rect 415400 148384 415452 148436
rect 99288 148316 99340 148368
rect 194784 148316 194836 148368
rect 370964 148316 371016 148368
rect 535460 148316 535512 148368
rect 156236 147636 156288 147688
rect 156420 147636 156472 147688
rect 168564 147636 168616 147688
rect 206008 147636 206060 147688
rect 226524 147636 226576 147688
rect 385132 147636 385184 147688
rect 385316 147636 385368 147688
rect 168656 147568 168708 147620
rect 206100 147568 206152 147620
rect 226616 147568 226668 147620
rect 324136 146956 324188 147008
rect 418160 146956 418212 147008
rect 103428 146888 103480 146940
rect 196072 146888 196124 146940
rect 373724 146888 373776 146940
rect 542360 146888 542412 146940
rect 107568 145528 107620 145580
rect 197544 145528 197596 145580
rect 353116 145528 353168 145580
rect 491300 145528 491352 145580
rect 181168 145027 181220 145036
rect 181168 144993 181177 145027
rect 181177 144993 181211 145027
rect 181211 144993 181220 145027
rect 181168 144984 181220 144993
rect 193496 144848 193548 144900
rect 193588 144848 193640 144900
rect 200304 144848 200356 144900
rect 200396 144848 200448 144900
rect 385224 144891 385276 144900
rect 385224 144857 385233 144891
rect 385233 144857 385267 144891
rect 385267 144857 385276 144891
rect 385224 144848 385276 144857
rect 110328 144168 110380 144220
rect 194140 144168 194192 144220
rect 358636 144168 358688 144220
rect 505100 144168 505152 144220
rect 158996 143531 159048 143540
rect 158996 143497 159005 143531
rect 159005 143497 159039 143531
rect 159039 143497 159048 143531
rect 158996 143488 159048 143497
rect 163228 143488 163280 143540
rect 168380 143488 168432 143540
rect 168656 143488 168708 143540
rect 179604 143531 179656 143540
rect 179604 143497 179613 143531
rect 179613 143497 179647 143531
rect 179647 143497 179656 143531
rect 179604 143488 179656 143497
rect 181168 143488 181220 143540
rect 183928 143488 183980 143540
rect 207296 143531 207348 143540
rect 207296 143497 207305 143531
rect 207305 143497 207339 143531
rect 207339 143497 207348 143531
rect 207296 143488 207348 143497
rect 219624 143531 219676 143540
rect 219624 143497 219633 143531
rect 219633 143497 219667 143531
rect 219667 143497 219676 143531
rect 219624 143488 219676 143497
rect 117228 142808 117280 142860
rect 201500 142808 201552 142860
rect 357256 142808 357308 142860
rect 502340 142808 502392 142860
rect 223856 142128 223908 142180
rect 121368 141380 121420 141432
rect 202972 141380 203024 141432
rect 355876 141380 355928 141432
rect 498200 141380 498252 141432
rect 125508 140020 125560 140072
rect 204536 140020 204588 140072
rect 362776 140020 362828 140072
rect 512092 140020 512144 140072
rect 46848 138660 46900 138712
rect 172612 138660 172664 138712
rect 361396 138660 361448 138712
rect 509240 138660 509292 138712
rect 240508 138116 240560 138168
rect 157616 138048 157668 138100
rect 217048 138048 217100 138100
rect 205916 137980 205968 138032
rect 206100 137980 206152 138032
rect 243084 138048 243136 138100
rect 242992 137980 243044 138032
rect 256884 137980 256936 138032
rect 157616 137912 157668 137964
rect 217048 137912 217100 137964
rect 256976 137912 257028 137964
rect 385224 137955 385276 137964
rect 385224 137921 385233 137955
rect 385233 137921 385267 137955
rect 385267 137921 385276 137955
rect 385224 137912 385276 137921
rect 57888 137232 57940 137284
rect 178224 137232 178276 137284
rect 341984 137232 342036 137284
rect 462320 137232 462372 137284
rect 3332 136552 3384 136604
rect 152924 136552 152976 136604
rect 344744 135872 344796 135924
rect 469220 135872 469272 135924
rect 210148 135192 210200 135244
rect 256976 135192 257028 135244
rect 257160 135192 257212 135244
rect 393044 135192 393096 135244
rect 579896 135192 579948 135244
rect 62028 134512 62080 134564
rect 181076 134011 181128 134020
rect 181076 133977 181085 134011
rect 181085 133977 181119 134011
rect 181119 133977 181128 134011
rect 181076 133968 181128 133977
rect 219624 134011 219676 134020
rect 219624 133977 219633 134011
rect 219633 133977 219667 134011
rect 219667 133977 219676 134011
rect 219624 133968 219676 133977
rect 240416 133943 240468 133952
rect 240416 133909 240425 133943
rect 240425 133909 240459 133943
rect 240459 133909 240468 133943
rect 240416 133900 240468 133909
rect 157800 133832 157852 133884
rect 181076 133875 181128 133884
rect 181076 133841 181085 133875
rect 181085 133841 181119 133875
rect 181119 133841 181128 133875
rect 181076 133832 181128 133841
rect 219624 133832 219676 133884
rect 219716 133832 219768 133884
rect 222476 133832 222528 133884
rect 343456 133152 343508 133204
rect 466460 133152 466512 133204
rect 378140 132472 378192 132524
rect 378324 132472 378376 132524
rect 347504 131724 347556 131776
rect 477592 131724 477644 131776
rect 159088 130976 159140 131028
rect 346216 130364 346268 130416
rect 473360 130364 473412 130416
rect 354496 129004 354548 129056
rect 492680 129004 492732 129056
rect 156236 128324 156288 128376
rect 156420 128324 156472 128376
rect 174084 128324 174136 128376
rect 174268 128324 174320 128376
rect 193404 128324 193456 128376
rect 193588 128324 193640 128376
rect 205732 128324 205784 128376
rect 205916 128324 205968 128376
rect 239036 128324 239088 128376
rect 163136 128299 163188 128308
rect 163136 128265 163145 128299
rect 163145 128265 163179 128299
rect 163179 128265 163188 128299
rect 163136 128256 163188 128265
rect 207296 128299 207348 128308
rect 207296 128265 207305 128299
rect 207305 128265 207339 128299
rect 207339 128265 207348 128299
rect 207296 128256 207348 128265
rect 210056 128299 210108 128308
rect 210056 128265 210065 128299
rect 210065 128265 210099 128299
rect 210099 128265 210108 128299
rect 210056 128256 210108 128265
rect 239128 128256 239180 128308
rect 348976 127576 349028 127628
rect 480260 127576 480312 127628
rect 372436 126216 372488 126268
rect 538220 126216 538272 126268
rect 182364 125536 182416 125588
rect 182456 125536 182508 125588
rect 196164 125579 196216 125588
rect 196164 125545 196173 125579
rect 196173 125545 196207 125579
rect 196207 125545 196216 125579
rect 196164 125536 196216 125545
rect 197636 125579 197688 125588
rect 197636 125545 197645 125579
rect 197645 125545 197679 125579
rect 197679 125545 197688 125579
rect 197636 125536 197688 125545
rect 216956 125536 217008 125588
rect 217048 125536 217100 125588
rect 218244 125536 218296 125588
rect 218428 125536 218480 125588
rect 221004 125536 221056 125588
rect 221188 125536 221240 125588
rect 364156 124856 364208 124908
rect 517520 124856 517572 124908
rect 183928 124244 183980 124296
rect 223856 124244 223908 124296
rect 157616 124219 157668 124228
rect 157616 124185 157625 124219
rect 157625 124185 157659 124219
rect 157659 124185 157668 124219
rect 157616 124176 157668 124185
rect 181168 124176 181220 124228
rect 222384 124219 222436 124228
rect 222384 124185 222393 124219
rect 222393 124185 222427 124219
rect 222427 124185 222436 124219
rect 222384 124176 222436 124185
rect 385040 124176 385092 124228
rect 385316 124176 385368 124228
rect 240416 124151 240468 124160
rect 240416 124117 240425 124151
rect 240425 124117 240459 124151
rect 240459 124117 240468 124151
rect 240416 124108 240468 124117
rect 392952 124108 393004 124160
rect 579896 124108 579948 124160
rect 223764 122859 223816 122868
rect 223764 122825 223773 122859
rect 223773 122825 223807 122859
rect 223807 122825 223816 122859
rect 223764 122816 223816 122825
rect 3332 122748 3384 122800
rect 153016 122748 153068 122800
rect 159088 122748 159140 122800
rect 183836 122748 183888 122800
rect 238760 122748 238812 122800
rect 239128 122748 239180 122800
rect 218428 119348 218480 119400
rect 219716 119348 219768 119400
rect 385040 119391 385092 119400
rect 385040 119357 385049 119391
rect 385049 119357 385083 119391
rect 385083 119357 385092 119391
rect 385040 119348 385092 119357
rect 163044 118668 163096 118720
rect 163228 118668 163280 118720
rect 174176 118668 174228 118720
rect 205824 118668 205876 118720
rect 207296 118668 207348 118720
rect 226616 118668 226668 118720
rect 256884 118668 256936 118720
rect 174268 118600 174320 118652
rect 205916 118600 205968 118652
rect 207388 118600 207440 118652
rect 226708 118600 226760 118652
rect 256976 118600 257028 118652
rect 181168 115991 181220 116000
rect 181168 115957 181177 115991
rect 181177 115957 181211 115991
rect 181211 115957 181220 115991
rect 181168 115948 181220 115957
rect 185124 115948 185176 116000
rect 185216 115948 185268 116000
rect 196164 115991 196216 116000
rect 196164 115957 196173 115991
rect 196173 115957 196207 115991
rect 196207 115957 196216 115991
rect 196164 115948 196216 115957
rect 197636 115991 197688 116000
rect 197636 115957 197645 115991
rect 197645 115957 197679 115991
rect 197679 115957 197688 115991
rect 197636 115948 197688 115957
rect 223764 115948 223816 116000
rect 225236 115948 225288 116000
rect 163136 115923 163188 115932
rect 163136 115889 163145 115923
rect 163145 115889 163179 115923
rect 163179 115889 163188 115923
rect 163136 115880 163188 115889
rect 222384 115880 222436 115932
rect 222568 115880 222620 115932
rect 223856 115812 223908 115864
rect 228088 115923 228140 115932
rect 228088 115889 228097 115923
rect 228097 115889 228131 115923
rect 228131 115889 228140 115923
rect 228088 115880 228140 115889
rect 256976 115880 257028 115932
rect 257160 115880 257212 115932
rect 225328 115812 225380 115864
rect 168564 114520 168616 114572
rect 168656 114520 168708 114572
rect 180984 114520 181036 114572
rect 218336 114563 218388 114572
rect 218336 114529 218345 114563
rect 218345 114529 218379 114563
rect 218379 114529 218388 114563
rect 218336 114520 218388 114529
rect 219624 114563 219676 114572
rect 219624 114529 219633 114563
rect 219633 114529 219667 114563
rect 219667 114529 219676 114563
rect 219624 114520 219676 114529
rect 240416 114563 240468 114572
rect 240416 114529 240425 114563
rect 240425 114529 240459 114563
rect 240459 114529 240468 114563
rect 240416 114520 240468 114529
rect 185124 114495 185176 114504
rect 185124 114461 185133 114495
rect 185133 114461 185167 114495
rect 185167 114461 185176 114495
rect 185124 114452 185176 114461
rect 180984 114427 181036 114436
rect 180984 114393 180993 114427
rect 180993 114393 181027 114427
rect 181027 114393 181036 114427
rect 180984 114384 181036 114393
rect 158904 113203 158956 113212
rect 158904 113169 158913 113203
rect 158913 113169 158947 113203
rect 158947 113169 158956 113203
rect 158904 113160 158956 113169
rect 183928 113203 183980 113212
rect 183928 113169 183937 113203
rect 183937 113169 183971 113203
rect 183971 113169 183980 113203
rect 183928 113160 183980 113169
rect 378140 113160 378192 113212
rect 378324 113160 378376 113212
rect 158904 113067 158956 113076
rect 158904 113033 158913 113067
rect 158913 113033 158947 113067
rect 158947 113033 158956 113067
rect 158904 113024 158956 113033
rect 395344 111732 395396 111784
rect 580172 111732 580224 111784
rect 225328 111188 225380 111240
rect 225236 111120 225288 111172
rect 185216 110984 185268 111036
rect 156236 109012 156288 109064
rect 156420 109012 156472 109064
rect 157616 109012 157668 109064
rect 174084 109012 174136 109064
rect 174268 109012 174320 109064
rect 193404 109012 193456 109064
rect 193588 109012 193640 109064
rect 205732 109012 205784 109064
rect 205916 109012 205968 109064
rect 157708 108944 157760 108996
rect 163136 108987 163188 108996
rect 163136 108953 163145 108987
rect 163145 108953 163179 108987
rect 163179 108953 163188 108987
rect 163136 108944 163188 108953
rect 218336 106292 218388 106344
rect 221096 106292 221148 106344
rect 228088 106335 228140 106344
rect 228088 106301 228097 106335
rect 228097 106301 228131 106335
rect 228131 106301 228140 106335
rect 228088 106292 228140 106301
rect 385040 106335 385092 106344
rect 385040 106301 385049 106335
rect 385049 106301 385083 106335
rect 385083 106301 385092 106335
rect 385040 106292 385092 106301
rect 196164 106267 196216 106276
rect 196164 106233 196173 106267
rect 196173 106233 196207 106267
rect 196207 106233 196216 106267
rect 196164 106224 196216 106233
rect 197636 106267 197688 106276
rect 197636 106233 197645 106267
rect 197645 106233 197679 106267
rect 197679 106233 197688 106267
rect 197636 106224 197688 106233
rect 200304 106224 200356 106276
rect 218244 106224 218296 106276
rect 221004 106224 221056 106276
rect 222568 106224 222620 106276
rect 238760 106224 238812 106276
rect 239036 106224 239088 106276
rect 240416 106267 240468 106276
rect 240416 106233 240425 106267
rect 240425 106233 240459 106267
rect 240459 106233 240468 106267
rect 240416 106224 240468 106233
rect 200304 106088 200356 106140
rect 219624 104932 219676 104984
rect 181168 104864 181220 104916
rect 182456 104907 182508 104916
rect 182456 104873 182465 104907
rect 182465 104873 182499 104907
rect 182499 104873 182508 104907
rect 182456 104864 182508 104873
rect 183836 104864 183888 104916
rect 183928 104864 183980 104916
rect 174176 104839 174228 104848
rect 174176 104805 174185 104839
rect 174185 104805 174219 104839
rect 174219 104805 174228 104839
rect 174176 104796 174228 104805
rect 385040 104839 385092 104848
rect 385040 104805 385049 104839
rect 385049 104805 385083 104839
rect 385083 104805 385092 104839
rect 385040 104796 385092 104805
rect 218244 104771 218296 104780
rect 218244 104737 218253 104771
rect 218253 104737 218287 104771
rect 218287 104737 218296 104771
rect 218244 104728 218296 104737
rect 219624 104728 219676 104780
rect 182364 103572 182416 103624
rect 159088 103504 159140 103556
rect 223856 103504 223908 103556
rect 223948 103368 224000 103420
rect 182456 102076 182508 102128
rect 183836 101396 183888 101448
rect 239036 101396 239088 101448
rect 183836 101260 183888 101312
rect 239036 101260 239088 101312
rect 218244 100011 218296 100020
rect 218244 99977 218253 100011
rect 218253 99977 218287 100011
rect 218287 99977 218296 100011
rect 218244 99968 218296 99977
rect 217048 99467 217100 99476
rect 217048 99433 217057 99467
rect 217057 99433 217091 99467
rect 217091 99433 217100 99467
rect 217048 99424 217100 99433
rect 157524 99356 157576 99408
rect 157708 99356 157760 99408
rect 163044 99356 163096 99408
rect 163228 99356 163280 99408
rect 181076 99356 181128 99408
rect 205824 99356 205876 99408
rect 207296 99356 207348 99408
rect 181168 99288 181220 99340
rect 205916 99288 205968 99340
rect 207388 99288 207440 99340
rect 219624 98676 219676 98728
rect 256700 97928 256752 97980
rect 256884 97928 256936 97980
rect 182456 97248 182508 97300
rect 196164 96679 196216 96688
rect 196164 96645 196173 96679
rect 196173 96645 196207 96679
rect 196207 96645 196216 96679
rect 196164 96636 196216 96645
rect 197636 96679 197688 96688
rect 197636 96645 197645 96679
rect 197645 96645 197679 96679
rect 197679 96645 197688 96679
rect 197636 96636 197688 96645
rect 222476 96679 222528 96688
rect 222476 96645 222485 96679
rect 222485 96645 222519 96679
rect 222519 96645 222528 96679
rect 222476 96636 222528 96645
rect 240416 96679 240468 96688
rect 240416 96645 240425 96679
rect 240425 96645 240459 96679
rect 240459 96645 240468 96679
rect 240416 96636 240468 96645
rect 163136 96611 163188 96620
rect 163136 96577 163145 96611
rect 163145 96577 163179 96611
rect 163179 96577 163188 96611
rect 163136 96568 163188 96577
rect 185032 96568 185084 96620
rect 185216 96568 185268 96620
rect 217048 96611 217100 96620
rect 217048 96577 217057 96611
rect 217057 96577 217091 96611
rect 217091 96577 217100 96611
rect 217048 96568 217100 96577
rect 158904 95208 158956 95260
rect 159088 95208 159140 95260
rect 168564 95208 168616 95260
rect 168656 95208 168708 95260
rect 174268 95208 174320 95260
rect 181076 95183 181128 95192
rect 181076 95149 181085 95183
rect 181085 95149 181119 95183
rect 181119 95149 181128 95183
rect 181076 95140 181128 95149
rect 185032 95183 185084 95192
rect 185032 95149 185041 95183
rect 185041 95149 185075 95183
rect 185075 95149 185084 95183
rect 185032 95140 185084 95149
rect 218244 95183 218296 95192
rect 218244 95149 218253 95183
rect 218253 95149 218287 95183
rect 218287 95149 218296 95183
rect 218244 95140 218296 95149
rect 158904 95115 158956 95124
rect 158904 95081 158913 95115
rect 158913 95081 158947 95115
rect 158947 95081 158956 95115
rect 158904 95072 158956 95081
rect 378140 93848 378192 93900
rect 378324 93848 378376 93900
rect 385132 93848 385184 93900
rect 3608 93780 3660 93832
rect 152740 93780 152792 93832
rect 227996 92463 228048 92472
rect 227996 92429 228005 92463
rect 228005 92429 228039 92463
rect 228039 92429 228048 92463
rect 227996 92420 228048 92429
rect 218336 91808 218388 91860
rect 156236 89700 156288 89752
rect 156420 89700 156472 89752
rect 157616 89700 157668 89752
rect 174084 89700 174136 89752
rect 174268 89700 174320 89752
rect 193404 89700 193456 89752
rect 193588 89700 193640 89752
rect 205732 89700 205784 89752
rect 205916 89700 205968 89752
rect 163136 89675 163188 89684
rect 163136 89641 163145 89675
rect 163145 89641 163179 89675
rect 163179 89641 163188 89675
rect 163136 89632 163188 89641
rect 157708 89564 157760 89616
rect 392860 88272 392912 88324
rect 579896 88272 579948 88324
rect 200304 86912 200356 86964
rect 209964 86912 210016 86964
rect 216956 86912 217008 86964
rect 217048 86912 217100 86964
rect 239036 86955 239088 86964
rect 239036 86921 239045 86955
rect 239045 86921 239079 86955
rect 239079 86921 239088 86955
rect 239036 86912 239088 86921
rect 240416 86955 240468 86964
rect 240416 86921 240425 86955
rect 240425 86921 240459 86955
rect 240459 86921 240468 86955
rect 240416 86912 240468 86921
rect 200304 86776 200356 86828
rect 183836 85799 183888 85808
rect 183836 85765 183845 85799
rect 183845 85765 183879 85799
rect 183879 85765 183888 85799
rect 183836 85756 183888 85765
rect 158996 85552 159048 85604
rect 181168 85552 181220 85604
rect 185216 85552 185268 85604
rect 221004 85552 221056 85604
rect 221096 85552 221148 85604
rect 223856 85552 223908 85604
rect 223948 85552 224000 85604
rect 174176 85527 174228 85536
rect 174176 85493 174185 85527
rect 174185 85493 174219 85527
rect 174219 85493 174228 85527
rect 174176 85484 174228 85493
rect 183836 84235 183888 84244
rect 183836 84201 183845 84235
rect 183845 84201 183879 84235
rect 183879 84201 183888 84235
rect 183836 84192 183888 84201
rect 182456 84167 182508 84176
rect 182456 84133 182465 84167
rect 182465 84133 182499 84167
rect 182499 84133 182508 84167
rect 182456 84124 182508 84133
rect 385132 84124 385184 84176
rect 228088 82832 228140 82884
rect 157524 80044 157576 80096
rect 157708 80044 157760 80096
rect 163044 80044 163096 80096
rect 163228 80044 163280 80096
rect 181076 80044 181128 80096
rect 205824 80044 205876 80096
rect 3056 79976 3108 80028
rect 152832 79976 152884 80028
rect 181168 79976 181220 80028
rect 207204 80112 207256 80164
rect 256884 80044 256936 80096
rect 207112 79976 207164 80028
rect 205916 79908 205968 79960
rect 256976 79908 257028 79960
rect 182456 79339 182508 79348
rect 182456 79305 182465 79339
rect 182465 79305 182499 79339
rect 182499 79305 182508 79339
rect 182456 79296 182508 79305
rect 228088 77936 228140 77988
rect 222568 77324 222620 77376
rect 209872 77299 209924 77308
rect 209872 77265 209881 77299
rect 209881 77265 209915 77299
rect 209915 77265 209924 77299
rect 209872 77256 209924 77265
rect 222476 77256 222528 77308
rect 239036 77299 239088 77308
rect 239036 77265 239045 77299
rect 239045 77265 239079 77299
rect 239079 77265 239088 77299
rect 239036 77256 239088 77265
rect 240416 77299 240468 77308
rect 240416 77265 240425 77299
rect 240425 77265 240459 77299
rect 240459 77265 240468 77299
rect 240416 77256 240468 77265
rect 207112 77231 207164 77240
rect 207112 77197 207121 77231
rect 207121 77197 207155 77231
rect 207155 77197 207164 77231
rect 207112 77188 207164 77197
rect 256976 77188 257028 77240
rect 392768 77188 392820 77240
rect 579896 77188 579948 77240
rect 158720 75896 158772 75948
rect 158904 75896 158956 75948
rect 174268 75896 174320 75948
rect 218244 75896 218296 75948
rect 218336 75896 218388 75948
rect 219624 75939 219676 75948
rect 219624 75905 219633 75939
rect 219633 75905 219667 75939
rect 219667 75905 219676 75939
rect 219624 75896 219676 75905
rect 181076 75871 181128 75880
rect 181076 75837 181085 75871
rect 181085 75837 181119 75871
rect 181119 75837 181128 75871
rect 181076 75828 181128 75837
rect 378140 74536 378192 74588
rect 378324 74536 378376 74588
rect 222476 73151 222528 73160
rect 222476 73117 222485 73151
rect 222485 73117 222519 73151
rect 222519 73117 222528 73151
rect 222476 73108 222528 73117
rect 183836 70703 183888 70712
rect 183836 70669 183845 70703
rect 183845 70669 183879 70703
rect 183879 70669 183888 70703
rect 183836 70660 183888 70669
rect 157616 70388 157668 70440
rect 163136 70388 163188 70440
rect 185124 70388 185176 70440
rect 157708 70252 157760 70304
rect 163228 70252 163280 70304
rect 207204 70320 207256 70372
rect 185216 70252 185268 70304
rect 205916 67668 205968 67720
rect 168564 67600 168616 67652
rect 168656 67600 168708 67652
rect 205824 67600 205876 67652
rect 256884 67643 256936 67652
rect 256884 67609 256893 67643
rect 256893 67609 256927 67643
rect 256927 67609 256936 67643
rect 256884 67600 256936 67609
rect 217048 67532 217100 67584
rect 240416 67575 240468 67584
rect 240416 67541 240425 67575
rect 240425 67541 240459 67575
rect 240459 67541 240468 67575
rect 240416 67532 240468 67541
rect 221096 66308 221148 66360
rect 225328 66308 225380 66360
rect 226708 66308 226760 66360
rect 174176 66240 174228 66292
rect 174268 66240 174320 66292
rect 181168 66240 181220 66292
rect 182364 66240 182416 66292
rect 182456 66240 182508 66292
rect 183836 66283 183888 66292
rect 183836 66249 183845 66283
rect 183845 66249 183879 66283
rect 183879 66249 183888 66283
rect 183836 66240 183888 66249
rect 221004 66240 221056 66292
rect 225236 66240 225288 66292
rect 226616 66240 226668 66292
rect 385040 66283 385092 66292
rect 385040 66249 385049 66283
rect 385049 66249 385083 66283
rect 385083 66249 385092 66283
rect 385040 66240 385092 66249
rect 158996 66215 159048 66224
rect 158996 66181 159005 66215
rect 159005 66181 159039 66215
rect 159039 66181 159048 66215
rect 158996 66172 159048 66181
rect 237288 66215 237340 66224
rect 237288 66181 237297 66215
rect 237297 66181 237331 66215
rect 237331 66181 237340 66215
rect 237288 66172 237340 66181
rect 238668 66215 238720 66224
rect 238668 66181 238677 66215
rect 238677 66181 238711 66215
rect 238711 66181 238720 66215
rect 238668 66172 238720 66181
rect 223764 64880 223816 64932
rect 223856 64880 223908 64932
rect 227996 64923 228048 64932
rect 227996 64889 228005 64923
rect 228005 64889 228039 64923
rect 228039 64889 228048 64923
rect 227996 64880 228048 64889
rect 182364 64855 182416 64864
rect 182364 64821 182373 64855
rect 182373 64821 182407 64855
rect 182407 64821 182416 64855
rect 182364 64812 182416 64821
rect 183836 64855 183888 64864
rect 183836 64821 183845 64855
rect 183845 64821 183879 64855
rect 183879 64821 183888 64855
rect 183836 64812 183888 64821
rect 185216 64855 185268 64864
rect 185216 64821 185225 64855
rect 185225 64821 185259 64855
rect 185259 64821 185268 64855
rect 185216 64812 185268 64821
rect 393964 64812 394016 64864
rect 580172 64812 580224 64864
rect 222660 63520 222712 63572
rect 240416 62747 240468 62756
rect 240416 62713 240425 62747
rect 240425 62713 240459 62747
rect 240459 62713 240468 62747
rect 240416 62704 240468 62713
rect 181168 60800 181220 60852
rect 207204 60664 207256 60716
rect 207388 60664 207440 60716
rect 209964 60664 210016 60716
rect 210148 60664 210200 60716
rect 185124 59168 185176 59220
rect 223764 58012 223816 58064
rect 168564 57944 168616 57996
rect 168656 57944 168708 57996
rect 219532 57944 219584 57996
rect 219624 57944 219676 57996
rect 221004 57944 221056 57996
rect 221096 57944 221148 57996
rect 225236 57944 225288 57996
rect 225328 57944 225380 57996
rect 256700 57944 256752 57996
rect 256976 57944 257028 57996
rect 180984 57919 181036 57928
rect 180984 57885 180993 57919
rect 180993 57885 181027 57919
rect 181027 57885 181036 57919
rect 180984 57876 181036 57885
rect 193588 57876 193640 57928
rect 210148 57876 210200 57928
rect 223764 57876 223816 57928
rect 239036 57919 239088 57928
rect 239036 57885 239045 57919
rect 239045 57885 239079 57919
rect 239079 57885 239088 57919
rect 239036 57876 239088 57885
rect 158996 56627 159048 56636
rect 158996 56593 159005 56627
rect 159005 56593 159039 56627
rect 159039 56593 159048 56627
rect 158996 56584 159048 56593
rect 217048 56584 217100 56636
rect 237288 56627 237340 56636
rect 237288 56593 237297 56627
rect 237297 56593 237331 56627
rect 237331 56593 237340 56627
rect 237288 56584 237340 56593
rect 238668 56627 238720 56636
rect 238668 56593 238677 56627
rect 238677 56593 238711 56627
rect 238711 56593 238720 56627
rect 238668 56584 238720 56593
rect 180984 56559 181036 56568
rect 180984 56525 180993 56559
rect 180993 56525 181027 56559
rect 181027 56525 181036 56559
rect 180984 56516 181036 56525
rect 218336 56516 218388 56568
rect 183836 55267 183888 55276
rect 183836 55233 183845 55267
rect 183845 55233 183879 55267
rect 183879 55233 183888 55267
rect 183836 55224 183888 55233
rect 378140 55224 378192 55276
rect 378324 55224 378376 55276
rect 222660 54612 222712 54664
rect 207388 51076 207440 51128
rect 3056 51008 3108 51060
rect 152556 51008 152608 51060
rect 207296 51008 207348 51060
rect 385132 51008 385184 51060
rect 385316 51008 385368 51060
rect 205916 48356 205968 48408
rect 219624 48356 219676 48408
rect 221096 48356 221148 48408
rect 158996 48288 159048 48340
rect 182364 48331 182416 48340
rect 182364 48297 182373 48331
rect 182373 48297 182407 48331
rect 182407 48297 182416 48331
rect 182364 48288 182416 48297
rect 193496 48331 193548 48340
rect 193496 48297 193505 48331
rect 193505 48297 193539 48331
rect 193539 48297 193548 48331
rect 193496 48288 193548 48297
rect 205824 48288 205876 48340
rect 210056 48331 210108 48340
rect 210056 48297 210065 48331
rect 210065 48297 210099 48331
rect 210099 48297 210108 48331
rect 210056 48288 210108 48297
rect 219532 48288 219584 48340
rect 221004 48288 221056 48340
rect 237196 48288 237248 48340
rect 237288 48288 237340 48340
rect 238668 48288 238720 48340
rect 238760 48288 238812 48340
rect 239036 48331 239088 48340
rect 239036 48297 239045 48331
rect 239045 48297 239079 48331
rect 239079 48297 239088 48331
rect 239036 48288 239088 48297
rect 256516 48288 256568 48340
rect 256884 48288 256936 48340
rect 158904 48220 158956 48272
rect 223764 48220 223816 48272
rect 223948 48220 224000 48272
rect 225236 48220 225288 48272
rect 225420 48220 225472 48272
rect 181168 46928 181220 46980
rect 218244 46971 218296 46980
rect 218244 46937 218253 46971
rect 218253 46937 218287 46971
rect 218287 46937 218296 46971
rect 218244 46928 218296 46937
rect 158904 46903 158956 46912
rect 158904 46869 158913 46903
rect 158913 46869 158947 46903
rect 158947 46869 158956 46903
rect 158904 46860 158956 46869
rect 182364 46903 182416 46912
rect 182364 46869 182373 46903
rect 182373 46869 182407 46903
rect 182407 46869 182416 46903
rect 182364 46860 182416 46869
rect 210056 46903 210108 46912
rect 210056 46869 210065 46903
rect 210065 46869 210099 46903
rect 210099 46869 210108 46903
rect 210056 46860 210108 46869
rect 221004 46903 221056 46912
rect 221004 46869 221013 46903
rect 221013 46869 221047 46903
rect 221047 46869 221056 46903
rect 221004 46860 221056 46869
rect 226616 46860 226668 46912
rect 226708 46860 226760 46912
rect 237288 46903 237340 46912
rect 237288 46869 237297 46903
rect 237297 46869 237331 46903
rect 237331 46869 237340 46903
rect 237288 46860 237340 46869
rect 238668 46903 238720 46912
rect 238668 46869 238677 46903
rect 238677 46869 238711 46903
rect 238711 46869 238720 46903
rect 238668 46860 238720 46869
rect 183928 45568 183980 45620
rect 184020 45568 184072 45620
rect 222568 45611 222620 45620
rect 222568 45577 222577 45611
rect 222577 45577 222611 45611
rect 222611 45577 222620 45611
rect 222568 45568 222620 45577
rect 185124 45500 185176 45552
rect 185400 45500 185452 45552
rect 181168 41420 181220 41472
rect 181076 41352 181128 41404
rect 392676 41352 392728 41404
rect 579896 41352 579948 41404
rect 219532 38743 219584 38752
rect 219532 38709 219541 38743
rect 219541 38709 219575 38743
rect 219575 38709 219584 38743
rect 219532 38700 219584 38709
rect 239036 38743 239088 38752
rect 239036 38709 239045 38743
rect 239045 38709 239079 38743
rect 239079 38709 239088 38743
rect 239036 38700 239088 38709
rect 168564 38632 168616 38684
rect 168656 38632 168708 38684
rect 218244 38632 218296 38684
rect 218336 38632 218388 38684
rect 256700 38632 256752 38684
rect 256976 38632 257028 38684
rect 163136 38607 163188 38616
rect 163136 38573 163145 38607
rect 163145 38573 163179 38607
rect 163179 38573 163188 38607
rect 163136 38564 163188 38573
rect 385408 38564 385460 38616
rect 182364 37315 182416 37324
rect 182364 37281 182373 37315
rect 182373 37281 182407 37315
rect 182407 37281 182416 37315
rect 182364 37272 182416 37281
rect 210148 37272 210200 37324
rect 221004 37315 221056 37324
rect 221004 37281 221013 37315
rect 221013 37281 221047 37315
rect 221047 37281 221056 37315
rect 221004 37272 221056 37281
rect 237288 37315 237340 37324
rect 237288 37281 237297 37315
rect 237297 37281 237331 37315
rect 237331 37281 237340 37315
rect 237288 37272 237340 37281
rect 238668 37315 238720 37324
rect 238668 37281 238677 37315
rect 238677 37281 238711 37315
rect 238711 37281 238720 37315
rect 238668 37272 238720 37281
rect 239036 37315 239088 37324
rect 239036 37281 239045 37315
rect 239045 37281 239079 37315
rect 239079 37281 239088 37315
rect 239036 37272 239088 37281
rect 207388 37247 207440 37256
rect 207388 37213 207397 37247
rect 207397 37213 207431 37247
rect 207431 37213 207440 37247
rect 207388 37204 207440 37213
rect 219532 35955 219584 35964
rect 219532 35921 219541 35955
rect 219541 35921 219575 35955
rect 219575 35921 219584 35955
rect 219532 35912 219584 35921
rect 378140 35912 378192 35964
rect 378324 35912 378376 35964
rect 3516 35844 3568 35896
rect 152648 35844 152700 35896
rect 181076 34731 181128 34740
rect 181076 34697 181085 34731
rect 181085 34697 181119 34731
rect 181119 34697 181128 34731
rect 181076 34688 181128 34697
rect 182364 31739 182416 31748
rect 182364 31705 182373 31739
rect 182373 31705 182407 31739
rect 182407 31705 182416 31739
rect 182364 31696 182416 31705
rect 205732 31696 205784 31748
rect 205916 31696 205968 31748
rect 225144 30336 225196 30388
rect 225420 30336 225472 30388
rect 392584 30268 392636 30320
rect 579896 30268 579948 30320
rect 159916 29588 159968 29640
rect 218336 29588 218388 29640
rect 158904 29087 158956 29096
rect 158904 29053 158913 29087
rect 158913 29053 158947 29087
rect 158947 29053 158956 29087
rect 158904 29044 158956 29053
rect 174268 29044 174320 29096
rect 163228 28976 163280 29028
rect 174176 28976 174228 29028
rect 181168 28976 181220 29028
rect 182364 29019 182416 29028
rect 182364 28985 182373 29019
rect 182373 28985 182407 29019
rect 182407 28985 182416 29019
rect 182364 28976 182416 28985
rect 216956 28976 217008 29028
rect 217048 28976 217100 29028
rect 256516 28976 256568 29028
rect 256792 28976 256844 29028
rect 385316 29019 385368 29028
rect 385316 28985 385325 29019
rect 385325 28985 385359 29019
rect 385359 28985 385368 29019
rect 385316 28976 385368 28985
rect 222384 28908 222436 28960
rect 222568 28908 222620 28960
rect 226616 28951 226668 28960
rect 226616 28917 226625 28951
rect 226625 28917 226659 28951
rect 226659 28917 226668 28951
rect 226616 28908 226668 28917
rect 239036 28951 239088 28960
rect 239036 28917 239045 28951
rect 239045 28917 239079 28951
rect 239079 28917 239088 28951
rect 239036 28908 239088 28917
rect 183468 28228 183520 28280
rect 228088 28228 228140 28280
rect 183928 27684 183980 27736
rect 223948 27684 224000 27736
rect 207388 27659 207440 27668
rect 207388 27625 207397 27659
rect 207397 27625 207431 27659
rect 207431 27625 207440 27659
rect 207388 27616 207440 27625
rect 223856 27616 223908 27668
rect 158904 27591 158956 27600
rect 158904 27557 158913 27591
rect 158913 27557 158947 27591
rect 158947 27557 158956 27591
rect 158904 27548 158956 27557
rect 181168 27591 181220 27600
rect 181168 27557 181177 27591
rect 181177 27557 181211 27591
rect 181211 27557 181220 27591
rect 181168 27548 181220 27557
rect 217048 27548 217100 27600
rect 219532 27591 219584 27600
rect 219532 27557 219541 27591
rect 219541 27557 219575 27591
rect 219575 27557 219584 27591
rect 219532 27548 219584 27557
rect 237288 27548 237340 27600
rect 238668 27548 238720 27600
rect 186228 26868 186280 26920
rect 229284 26868 229336 26920
rect 183744 26367 183796 26376
rect 183744 26333 183753 26367
rect 183753 26333 183787 26367
rect 183787 26333 183796 26367
rect 183744 26324 183796 26333
rect 183744 26231 183796 26240
rect 183744 26197 183753 26231
rect 183753 26197 183787 26231
rect 183787 26197 183796 26231
rect 183744 26188 183796 26197
rect 157248 25508 157300 25560
rect 215944 25508 215996 25560
rect 153108 24080 153160 24132
rect 214564 24080 214616 24132
rect 141976 22720 142028 22772
rect 211252 22720 211304 22772
rect 239036 22763 239088 22772
rect 239036 22729 239045 22763
rect 239045 22729 239079 22763
rect 239079 22729 239088 22763
rect 239036 22720 239088 22729
rect 182364 22108 182416 22160
rect 207388 22108 207440 22160
rect 221096 22108 221148 22160
rect 156236 22040 156288 22092
rect 156420 22040 156472 22092
rect 200304 22040 200356 22092
rect 182456 21972 182508 22024
rect 256884 22040 256936 22092
rect 257068 22040 257120 22092
rect 200396 21972 200448 22024
rect 221096 21972 221148 22024
rect 188988 21360 189040 21412
rect 230664 21360 230716 21412
rect 292304 21360 292356 21412
rect 339592 21360 339644 21412
rect 365536 21360 365588 21412
rect 520372 21360 520424 21412
rect 180708 19932 180760 19984
rect 291016 19932 291068 19984
rect 336740 19932 336792 19984
rect 361488 19932 361540 19984
rect 510620 19932 510672 19984
rect 156420 19295 156472 19304
rect 156420 19261 156429 19295
rect 156429 19261 156463 19295
rect 156463 19261 156472 19295
rect 156420 19252 156472 19261
rect 200396 19295 200448 19304
rect 200396 19261 200405 19295
rect 200405 19261 200439 19295
rect 200439 19261 200448 19295
rect 200396 19252 200448 19261
rect 222476 19295 222528 19304
rect 222476 19261 222485 19295
rect 222485 19261 222519 19295
rect 222519 19261 222528 19295
rect 222476 19252 222528 19261
rect 257068 19295 257120 19304
rect 257068 19261 257077 19295
rect 257077 19261 257111 19295
rect 257111 19261 257120 19295
rect 257068 19252 257120 19261
rect 385132 19252 385184 19304
rect 158904 19227 158956 19236
rect 158904 19193 158913 19227
rect 158913 19193 158947 19227
rect 158947 19193 158956 19227
rect 158904 19184 158956 19193
rect 173808 18572 173860 18624
rect 223856 18572 223908 18624
rect 286784 18572 286836 18624
rect 325700 18572 325752 18624
rect 360108 18572 360160 18624
rect 506480 18572 506532 18624
rect 181168 18003 181220 18012
rect 181168 17969 181177 18003
rect 181177 17969 181211 18003
rect 181211 17969 181220 18003
rect 181168 17960 181220 17969
rect 185124 17960 185176 18012
rect 185400 17960 185452 18012
rect 207204 18003 207256 18012
rect 207204 17969 207213 18003
rect 207213 17969 207247 18003
rect 207247 17969 207256 18003
rect 207204 17960 207256 17969
rect 135168 17212 135220 17264
rect 208400 17212 208452 17264
rect 281356 17212 281408 17264
rect 311900 17212 311952 17264
rect 358728 17212 358780 17264
rect 502432 17212 502484 17264
rect 183744 16643 183796 16652
rect 183744 16609 183753 16643
rect 183753 16609 183787 16643
rect 183787 16609 183796 16643
rect 183744 16600 183796 16609
rect 378140 16600 378192 16652
rect 378324 16600 378376 16652
rect 187608 15852 187660 15904
rect 229192 15852 229244 15904
rect 277124 15852 277176 15904
rect 300860 15852 300912 15904
rect 357348 15852 357400 15904
rect 499580 15852 499632 15904
rect 180984 14492 181036 14544
rect 181168 14492 181220 14544
rect 184848 14424 184900 14476
rect 227812 14424 227864 14476
rect 285404 14424 285456 14476
rect 321652 14424 321704 14476
rect 354588 14424 354640 14476
rect 494152 14424 494204 14476
rect 183744 13175 183796 13184
rect 183744 13141 183753 13175
rect 183753 13141 183787 13175
rect 183787 13141 183796 13175
rect 183744 13132 183796 13141
rect 278596 13132 278648 13184
rect 305000 13132 305052 13184
rect 176568 13064 176620 13116
rect 225144 13064 225196 13116
rect 282644 13064 282696 13116
rect 314660 13064 314712 13116
rect 355968 13064 356020 13116
rect 495440 13064 495492 13116
rect 185124 12495 185176 12504
rect 185124 12461 185133 12495
rect 185133 12461 185167 12495
rect 185167 12461 185176 12495
rect 185124 12452 185176 12461
rect 156420 12427 156472 12436
rect 156420 12393 156429 12427
rect 156429 12393 156463 12427
rect 156463 12393 156472 12427
rect 156420 12384 156472 12393
rect 205732 12384 205784 12436
rect 205916 12384 205968 12436
rect 257068 12291 257120 12300
rect 257068 12257 257077 12291
rect 257077 12257 257111 12291
rect 257111 12257 257120 12291
rect 257068 12248 257120 12257
rect 279976 11772 280028 11824
rect 307760 11772 307812 11824
rect 23388 11704 23440 11756
rect 164332 11704 164384 11756
rect 169392 11704 169444 11756
rect 289544 11704 289596 11756
rect 332600 11704 332652 11756
rect 351736 11704 351788 11756
rect 485872 11704 485924 11756
rect 192024 10344 192076 10396
rect 231952 10344 232004 10396
rect 278688 10344 278740 10396
rect 305092 10344 305144 10396
rect 13636 10276 13688 10328
rect 160192 10276 160244 10328
rect 165896 10276 165948 10328
rect 221096 10276 221148 10328
rect 288256 10276 288308 10328
rect 329840 10276 329892 10328
rect 353208 10276 353260 10328
rect 488540 10276 488592 10328
rect 158904 9664 158956 9716
rect 158996 9664 159048 9716
rect 200396 9707 200448 9716
rect 200396 9673 200405 9707
rect 200405 9673 200439 9707
rect 200439 9673 200448 9707
rect 200396 9664 200448 9673
rect 216956 9707 217008 9716
rect 216956 9673 216965 9707
rect 216965 9673 216999 9707
rect 216999 9673 217008 9707
rect 216956 9664 217008 9673
rect 219532 9707 219584 9716
rect 219532 9673 219541 9707
rect 219541 9673 219575 9707
rect 219575 9673 219584 9707
rect 219532 9664 219584 9673
rect 237196 9707 237248 9716
rect 237196 9673 237205 9707
rect 237205 9673 237239 9707
rect 237239 9673 237248 9707
rect 237196 9664 237248 9673
rect 238392 9707 238444 9716
rect 238392 9673 238401 9707
rect 238401 9673 238435 9707
rect 238435 9673 238444 9707
rect 238392 9664 238444 9673
rect 385040 9707 385092 9716
rect 385040 9673 385049 9707
rect 385049 9673 385083 9707
rect 385083 9673 385092 9707
rect 385040 9664 385092 9673
rect 312544 9596 312596 9648
rect 313372 9596 313424 9648
rect 326896 9596 326948 9648
rect 423956 9596 424008 9648
rect 328184 9528 328236 9580
rect 427544 9528 427596 9580
rect 329656 9460 329708 9512
rect 431132 9460 431184 9512
rect 330944 9392 330996 9444
rect 434628 9392 434680 9444
rect 332416 9324 332468 9376
rect 438216 9324 438268 9376
rect 333704 9256 333756 9308
rect 441804 9256 441856 9308
rect 335176 9188 335228 9240
rect 445392 9188 445444 9240
rect 336556 9120 336608 9172
rect 448980 9120 449032 9172
rect 337936 9052 337988 9104
rect 452476 9052 452528 9104
rect 184756 8984 184808 9036
rect 229100 8984 229152 9036
rect 278044 8984 278096 9036
rect 299112 8984 299164 9036
rect 339224 8984 339276 9036
rect 456064 8984 456116 9036
rect 162308 8916 162360 8968
rect 219532 8916 219584 8968
rect 275836 8916 275888 8968
rect 297732 8916 297784 8968
rect 340696 8916 340748 8968
rect 459652 8916 459704 8968
rect 324228 8848 324280 8900
rect 420368 8848 420420 8900
rect 322756 8780 322808 8832
rect 416872 8780 416924 8832
rect 321468 8712 321520 8764
rect 413284 8712 413336 8764
rect 319996 8644 320048 8696
rect 409696 8644 409748 8696
rect 318708 8576 318760 8628
rect 406108 8576 406160 8628
rect 317236 8508 317288 8560
rect 402520 8508 402572 8560
rect 315948 8440 316000 8492
rect 399024 8440 399076 8492
rect 3424 8236 3476 8288
rect 152464 8236 152516 8288
rect 375104 8236 375156 8288
rect 545304 8236 545356 8288
rect 94504 8168 94556 8220
rect 191932 8168 191984 8220
rect 299204 8168 299256 8220
rect 356152 8168 356204 8220
rect 376484 8168 376536 8220
rect 548892 8168 548944 8220
rect 77852 8100 77904 8152
rect 186504 8100 186556 8152
rect 300584 8100 300636 8152
rect 359740 8100 359792 8152
rect 377864 8100 377916 8152
rect 552388 8100 552440 8152
rect 74264 8032 74316 8084
rect 302056 8032 302108 8084
rect 363328 8032 363380 8084
rect 379244 8032 379296 8084
rect 555976 8032 556028 8084
rect 70676 7964 70728 8016
rect 182364 7964 182416 8016
rect 303344 7964 303396 8016
rect 366916 7964 366968 8016
rect 380624 7964 380676 8016
rect 559564 7964 559616 8016
rect 67180 7896 67232 7948
rect 180984 7896 181036 7948
rect 304724 7896 304776 7948
rect 370412 7896 370464 7948
rect 382004 7896 382056 7948
rect 563152 7896 563204 7948
rect 63592 7828 63644 7880
rect 179512 7828 179564 7880
rect 306104 7828 306156 7880
rect 374000 7828 374052 7880
rect 383476 7828 383528 7880
rect 566740 7828 566792 7880
rect 60004 7760 60056 7812
rect 178132 7760 178184 7812
rect 307576 7760 307628 7812
rect 377588 7760 377640 7812
rect 384764 7760 384816 7812
rect 570236 7760 570288 7812
rect 56416 7692 56468 7744
rect 176752 7692 176804 7744
rect 308864 7692 308916 7744
rect 381176 7692 381228 7744
rect 386144 7692 386196 7744
rect 573824 7692 573876 7744
rect 52828 7624 52880 7676
rect 175372 7624 175424 7676
rect 271604 7624 271656 7676
rect 287152 7624 287204 7676
rect 310336 7624 310388 7676
rect 384672 7624 384724 7676
rect 387524 7624 387576 7676
rect 577412 7624 577464 7676
rect 49332 7556 49384 7608
rect 174084 7556 174136 7608
rect 201500 7556 201552 7608
rect 236092 7556 236144 7608
rect 274456 7556 274508 7608
rect 295524 7556 295576 7608
rect 311624 7556 311676 7608
rect 388260 7556 388312 7608
rect 388904 7556 388956 7608
rect 581000 7556 581052 7608
rect 98092 7488 98144 7540
rect 193312 7488 193364 7540
rect 373816 7488 373868 7540
rect 541716 7488 541768 7540
rect 101588 7420 101640 7472
rect 194692 7420 194744 7472
rect 372528 7420 372580 7472
rect 538128 7420 538180 7472
rect 105176 7352 105228 7404
rect 197452 7352 197504 7404
rect 371056 7352 371108 7404
rect 534540 7352 534592 7404
rect 108764 7284 108816 7336
rect 198924 7284 198976 7336
rect 369676 7284 369728 7336
rect 531044 7284 531096 7336
rect 112352 7216 112404 7268
rect 200212 7216 200264 7268
rect 368296 7216 368348 7268
rect 527456 7216 527508 7268
rect 115940 7148 115992 7200
rect 201684 7148 201736 7200
rect 366824 7148 366876 7200
rect 523868 7148 523920 7200
rect 119436 7080 119488 7132
rect 203064 7080 203116 7132
rect 314476 7080 314528 7132
rect 395436 7080 395488 7132
rect 123024 7012 123076 7064
rect 204352 7012 204404 7064
rect 313188 7012 313240 7064
rect 391848 7012 391900 7064
rect 132592 6808 132644 6860
rect 207296 6808 207348 6860
rect 338028 6808 338080 6860
rect 451280 6808 451332 6860
rect 129004 6740 129056 6792
rect 205732 6740 205784 6792
rect 339316 6740 339368 6792
rect 454868 6740 454920 6792
rect 90916 6672 90968 6724
rect 190552 6672 190604 6724
rect 340788 6672 340840 6724
rect 458456 6672 458508 6724
rect 87328 6604 87380 6656
rect 189172 6604 189224 6656
rect 342076 6604 342128 6656
rect 462044 6604 462096 6656
rect 83832 6536 83884 6588
rect 187792 6536 187844 6588
rect 343548 6536 343600 6588
rect 465632 6536 465684 6588
rect 44548 6468 44600 6520
rect 172520 6468 172572 6520
rect 344836 6468 344888 6520
rect 469128 6468 469180 6520
rect 40960 6400 41012 6452
rect 171232 6400 171284 6452
rect 178960 6400 179012 6452
rect 226432 6400 226484 6452
rect 346308 6400 346360 6452
rect 472716 6400 472768 6452
rect 37372 6332 37424 6384
rect 169852 6332 169904 6384
rect 175372 6332 175424 6384
rect 225052 6332 225104 6384
rect 347596 6332 347648 6384
rect 476304 6332 476356 6384
rect 33876 6264 33928 6316
rect 168472 6264 168524 6316
rect 171784 6264 171836 6316
rect 223672 6264 223724 6316
rect 349068 6264 349120 6316
rect 479892 6264 479944 6316
rect 8852 6196 8904 6248
rect 157432 6196 157484 6248
rect 161112 6196 161164 6248
rect 219440 6196 219492 6248
rect 277216 6196 277268 6248
rect 302608 6196 302660 6248
rect 350356 6196 350408 6248
rect 484584 6196 484636 6248
rect 4068 6128 4120 6180
rect 156144 6128 156196 6180
rect 157524 6128 157576 6180
rect 218152 6128 218204 6180
rect 272984 6128 273036 6180
rect 136088 6060 136140 6112
rect 210056 6060 210108 6112
rect 139676 5992 139728 6044
rect 211344 5992 211396 6044
rect 290464 6128 290516 6180
rect 319260 6128 319312 6180
rect 351828 6128 351880 6180
rect 488172 6128 488224 6180
rect 335268 6060 335320 6112
rect 447784 6060 447836 6112
rect 290740 5992 290792 6044
rect 333796 5992 333848 6044
rect 444196 5992 444248 6044
rect 143264 5924 143316 5976
rect 212540 5924 212592 5976
rect 332508 5924 332560 5976
rect 440608 5924 440660 5976
rect 146852 5856 146904 5908
rect 213920 5856 213972 5908
rect 331036 5856 331088 5908
rect 437020 5856 437072 5908
rect 150440 5788 150492 5840
rect 215484 5788 215536 5840
rect 230480 5788 230532 5840
rect 329748 5788 329800 5840
rect 433524 5788 433576 5840
rect 153936 5720 153988 5772
rect 216772 5720 216824 5772
rect 328276 5720 328328 5772
rect 429936 5720 429988 5772
rect 164700 5652 164752 5704
rect 220912 5652 220964 5704
rect 326988 5652 327040 5704
rect 426348 5652 426400 5704
rect 168196 5584 168248 5636
rect 222292 5584 222344 5636
rect 325516 5584 325568 5636
rect 422760 5584 422812 5636
rect 287704 5516 287756 5568
rect 294328 5516 294380 5568
rect 51632 5448 51684 5500
rect 175280 5448 175332 5500
rect 198004 5448 198056 5500
rect 234712 5448 234764 5500
rect 296444 5448 296496 5500
rect 351368 5448 351420 5500
rect 375196 5448 375248 5500
rect 544108 5448 544160 5500
rect 48136 5380 48188 5432
rect 173992 5380 174044 5432
rect 190828 5380 190880 5432
rect 230572 5380 230624 5432
rect 297824 5380 297876 5432
rect 354956 5380 355008 5432
rect 376576 5380 376628 5432
rect 547696 5380 547748 5432
rect 30288 5312 30340 5364
rect 167184 5312 167236 5364
rect 194508 5312 194560 5364
rect 233332 5312 233384 5364
rect 299296 5312 299348 5364
rect 358544 5312 358596 5364
rect 377956 5312 378008 5364
rect 551192 5312 551244 5364
rect 26700 5244 26752 5296
rect 165712 5244 165764 5296
rect 181352 5244 181404 5296
rect 227720 5244 227772 5296
rect 300676 5244 300728 5296
rect 362132 5244 362184 5296
rect 379336 5244 379388 5296
rect 554780 5244 554832 5296
rect 21916 5176 21968 5228
rect 163136 5176 163188 5228
rect 177764 5176 177816 5228
rect 226340 5176 226392 5228
rect 303436 5176 303488 5228
rect 365720 5176 365772 5228
rect 380716 5176 380768 5228
rect 558368 5176 558420 5228
rect 17224 5108 17276 5160
rect 161480 5108 161532 5160
rect 174176 5108 174228 5160
rect 224960 5108 225012 5160
rect 304816 5108 304868 5160
rect 369216 5108 369268 5160
rect 382096 5108 382148 5160
rect 561956 5108 562008 5160
rect 12440 5040 12492 5092
rect 158812 5040 158864 5092
rect 170588 5040 170640 5092
rect 223580 5040 223632 5092
rect 306196 5040 306248 5092
rect 372804 5040 372856 5092
rect 383568 5040 383620 5092
rect 565544 5040 565596 5092
rect 7656 4972 7708 5024
rect 157708 4972 157760 5024
rect 167092 4972 167144 5024
rect 222200 4972 222252 5024
rect 307668 4972 307720 5024
rect 376392 4972 376444 5024
rect 384856 4972 384908 5024
rect 569040 4972 569092 5024
rect 1676 4904 1728 4956
rect 154580 4904 154632 4956
rect 163504 4904 163556 4956
rect 220820 4904 220872 4956
rect 308956 4904 309008 4956
rect 379980 4904 380032 4956
rect 386236 4904 386288 4956
rect 572628 4904 572680 4956
rect 2872 4836 2924 4888
rect 156052 4836 156104 4888
rect 158720 4836 158772 4888
rect 218060 4836 218112 4888
rect 310428 4836 310480 4888
rect 383568 4836 383620 4888
rect 387616 4836 387668 4888
rect 576216 4836 576268 4888
rect 572 4768 624 4820
rect 154672 4768 154724 4820
rect 155132 4768 155184 4820
rect 216956 4768 217008 4820
rect 233424 4768 233476 4820
rect 270224 4768 270276 4820
rect 283656 4768 283708 4820
rect 311716 4768 311768 4820
rect 387064 4768 387116 4820
rect 388996 4768 389048 4820
rect 579804 4768 579856 4820
rect 55220 4700 55272 4752
rect 176660 4700 176712 4752
rect 297916 4700 297968 4752
rect 352564 4700 352616 4752
rect 371148 4700 371200 4752
rect 536932 4700 536984 4752
rect 58808 4632 58860 4684
rect 178040 4632 178092 4684
rect 295156 4632 295208 4684
rect 347872 4632 347924 4684
rect 373908 4632 373960 4684
rect 540520 4632 540572 4684
rect 62396 4564 62448 4616
rect 179420 4564 179472 4616
rect 296536 4564 296588 4616
rect 349068 4564 349120 4616
rect 369768 4564 369820 4616
rect 533436 4564 533488 4616
rect 65984 4496 66036 4548
rect 180892 4496 180944 4548
rect 293684 4496 293736 4548
rect 344284 4496 344336 4548
rect 368388 4496 368440 4548
rect 529848 4496 529900 4548
rect 69480 4428 69532 4480
rect 182272 4428 182324 4480
rect 295064 4428 295116 4480
rect 345480 4428 345532 4480
rect 367008 4428 367060 4480
rect 526260 4428 526312 4480
rect 73068 4360 73120 4412
rect 183652 4360 183704 4412
rect 293776 4360 293828 4412
rect 341892 4360 341944 4412
rect 365628 4360 365680 4412
rect 522672 4360 522724 4412
rect 76656 4292 76708 4344
rect 292396 4292 292448 4344
rect 338304 4292 338356 4344
rect 364248 4292 364300 4344
rect 519084 4292 519136 4344
rect 80244 4224 80296 4276
rect 186412 4224 186464 4276
rect 289636 4224 289688 4276
rect 334716 4224 334768 4276
rect 362868 4224 362920 4276
rect 515588 4224 515640 4276
rect 140872 4156 140924 4208
rect 142068 4156 142120 4208
rect 14832 4088 14884 4140
rect 18604 4088 18656 4140
rect 187700 4088 187752 4140
rect 188436 4088 188488 4140
rect 188988 4088 189040 4140
rect 199200 4088 199252 4140
rect 200028 4088 200080 4140
rect 200396 4088 200448 4140
rect 201408 4088 201460 4140
rect 206284 4088 206336 4140
rect 206928 4088 206980 4140
rect 215852 4088 215904 4140
rect 216588 4088 216640 4140
rect 217048 4088 217100 4140
rect 217968 4088 218020 4140
rect 218152 4088 218204 4140
rect 222936 4088 222988 4140
rect 223488 4088 223540 4140
rect 234804 4088 234856 4140
rect 235908 4088 235960 4140
rect 240784 4088 240836 4140
rect 241428 4088 241480 4140
rect 82636 4020 82688 4072
rect 186320 4020 186372 4072
rect 221740 4020 221792 4072
rect 244280 4088 244332 4140
rect 244372 4088 244424 4140
rect 245568 4088 245620 4140
rect 257436 4088 257488 4140
rect 257988 4088 258040 4140
rect 258172 4088 258224 4140
rect 258632 4088 258684 4140
rect 262128 4088 262180 4140
rect 263416 4088 263468 4140
rect 270316 4088 270368 4140
rect 284760 4088 284812 4140
rect 289728 4088 289780 4140
rect 332416 4088 332468 4140
rect 339408 4088 339460 4140
rect 457260 4088 457312 4140
rect 243176 4020 243228 4072
rect 244924 4020 244976 4072
rect 260748 4020 260800 4072
rect 262220 4020 262272 4072
rect 270408 4020 270460 4072
rect 285956 4020 286008 4072
rect 291108 4020 291160 4072
rect 335912 4020 335964 4072
rect 342168 4020 342220 4072
rect 464436 4020 464488 4072
rect 75460 3952 75512 4004
rect 71872 3884 71924 3936
rect 68284 3816 68336 3868
rect 172980 3816 173032 3868
rect 173808 3816 173860 3868
rect 64788 3748 64840 3800
rect 180156 3952 180208 4004
rect 180708 3952 180760 4004
rect 182548 3952 182600 4004
rect 183468 3952 183520 4004
rect 208676 3952 208728 4004
rect 220544 3952 220596 4004
rect 241612 3952 241664 4004
rect 267004 3952 267056 4004
rect 270500 3952 270552 4004
rect 271696 3952 271748 4004
rect 288348 3952 288400 4004
rect 292488 3952 292540 4004
rect 339500 3952 339552 4004
rect 344928 3952 344980 4004
rect 471520 3952 471572 4004
rect 214656 3884 214708 3936
rect 226524 3884 226576 3936
rect 227628 3884 227680 3936
rect 184940 3816 184992 3868
rect 209872 3816 209924 3868
rect 183560 3748 183612 3800
rect 240232 3884 240284 3936
rect 264244 3884 264296 3936
rect 268108 3884 268160 3936
rect 271788 3884 271840 3936
rect 289544 3884 289596 3936
rect 293868 3884 293920 3936
rect 343088 3884 343140 3936
rect 347688 3884 347740 3936
rect 478696 3884 478748 3936
rect 485780 3884 485832 3936
rect 486976 3884 487028 3936
rect 494152 3884 494204 3936
rect 495348 3884 495400 3936
rect 502432 3884 502484 3936
rect 503628 3884 503680 3936
rect 239036 3816 239088 3868
rect 268844 3816 268896 3868
rect 46940 3680 46992 3732
rect 173900 3680 173952 3732
rect 180800 3680 180852 3732
rect 238852 3748 238904 3800
rect 264796 3748 264848 3800
rect 271696 3748 271748 3800
rect 230112 3680 230164 3732
rect 231124 3680 231176 3732
rect 233700 3680 233752 3732
rect 234528 3680 234580 3732
rect 242900 3680 242952 3732
rect 264888 3680 264940 3732
rect 272892 3680 272944 3732
rect 273076 3816 273128 3868
rect 291936 3816 291988 3868
rect 295248 3816 295300 3868
rect 346676 3816 346728 3868
rect 375288 3816 375340 3868
rect 546500 3816 546552 3868
rect 273168 3748 273220 3800
rect 293132 3748 293184 3800
rect 296628 3748 296680 3800
rect 350264 3748 350316 3800
rect 376668 3748 376720 3800
rect 550088 3748 550140 3800
rect 34980 3612 35032 3664
rect 36544 3612 36596 3664
rect 43352 3612 43404 3664
rect 165804 3612 165856 3664
rect 39764 3544 39816 3596
rect 169760 3544 169812 3596
rect 182180 3612 182232 3664
rect 193220 3612 193272 3664
rect 194416 3612 194468 3664
rect 207480 3612 207532 3664
rect 237472 3612 237524 3664
rect 240416 3544 240468 3596
rect 16028 3476 16080 3528
rect 19984 3476 20036 3528
rect 25504 3476 25556 3528
rect 29644 3476 29696 3528
rect 31484 3476 31536 3528
rect 32404 3476 32456 3528
rect 32680 3476 32732 3528
rect 35164 3476 35216 3528
rect 42156 3476 42208 3528
rect 42708 3476 42760 3528
rect 168748 3476 168800 3528
rect 183744 3476 183796 3528
rect 184848 3476 184900 3528
rect 237564 3476 237616 3528
rect 241980 3476 242032 3528
rect 242808 3476 242860 3528
rect 251364 3612 251416 3664
rect 266176 3612 266228 3664
rect 274088 3612 274140 3664
rect 274548 3680 274600 3732
rect 296720 3680 296772 3732
rect 298008 3680 298060 3732
rect 275928 3612 275980 3664
rect 300308 3612 300360 3664
rect 300768 3680 300820 3732
rect 305000 3680 305052 3732
rect 306104 3680 306156 3732
rect 353760 3680 353812 3732
rect 378048 3680 378100 3732
rect 553584 3680 553636 3732
rect 360936 3612 360988 3664
rect 379428 3612 379480 3664
rect 557172 3612 557224 3664
rect 266268 3544 266320 3596
rect 276480 3544 276532 3596
rect 277308 3544 277360 3596
rect 303804 3544 303856 3596
rect 304908 3544 304960 3596
rect 371608 3544 371660 3596
rect 380808 3544 380860 3596
rect 560760 3544 560812 3596
rect 6460 3408 6512 3460
rect 10324 3408 10376 3460
rect 29092 3408 29144 3460
rect 171140 3408 171192 3460
rect 189632 3408 189684 3460
rect 45744 3340 45796 3392
rect 46848 3340 46900 3392
rect 50528 3340 50580 3392
rect 50988 3340 51040 3392
rect 54024 3340 54076 3392
rect 55128 3340 55180 3392
rect 61200 3340 61252 3392
rect 62028 3340 62080 3392
rect 81440 3340 81492 3392
rect 82728 3340 82780 3392
rect 18328 3272 18380 3324
rect 21364 3272 21416 3324
rect 36176 3272 36228 3324
rect 27896 3204 27948 3256
rect 31024 3204 31076 3256
rect 79048 3204 79100 3256
rect 84936 3340 84988 3392
rect 85488 3340 85540 3392
rect 88524 3340 88576 3392
rect 89628 3340 89680 3392
rect 86132 3204 86184 3256
rect 189080 3340 189132 3392
rect 212264 3408 212316 3460
rect 239588 3408 239640 3460
rect 249156 3476 249208 3528
rect 249708 3476 249760 3528
rect 252652 3476 252704 3528
rect 253848 3476 253900 3528
rect 267648 3476 267700 3528
rect 277676 3476 277728 3528
rect 280068 3476 280120 3528
rect 307392 3476 307444 3528
rect 309048 3476 309100 3528
rect 382372 3476 382424 3528
rect 384948 3476 385000 3528
rect 567844 3476 567896 3528
rect 249892 3408 249944 3460
rect 267556 3408 267608 3460
rect 278872 3408 278924 3460
rect 281448 3408 281500 3460
rect 310980 3408 311032 3460
rect 311808 3408 311860 3460
rect 389456 3408 389508 3460
rect 390468 3408 390520 3460
rect 582196 3408 582248 3460
rect 89904 3272 89956 3324
rect 190736 3272 190788 3324
rect 225328 3340 225380 3392
rect 245752 3340 245804 3392
rect 269028 3340 269080 3392
rect 93308 3204 93360 3256
rect 192116 3204 192168 3256
rect 95700 3136 95752 3188
rect 96528 3136 96580 3188
rect 102784 3136 102836 3188
rect 103428 3136 103480 3188
rect 106372 3136 106424 3188
rect 107568 3136 107620 3188
rect 111156 3136 111208 3188
rect 111708 3136 111760 3188
rect 193404 3136 193456 3188
rect 100484 3068 100536 3120
rect 194600 3068 194652 3120
rect 96896 3000 96948 3052
rect 196164 3000 196216 3052
rect 196808 3000 196860 3052
rect 197268 3000 197320 3052
rect 227720 3272 227772 3324
rect 229008 3272 229060 3324
rect 228916 3204 228968 3256
rect 247132 3272 247184 3324
rect 268384 3272 268436 3324
rect 275284 3272 275336 3324
rect 282460 3340 282512 3392
rect 286876 3340 286928 3392
rect 327632 3340 327684 3392
rect 336648 3340 336700 3392
rect 450176 3340 450228 3392
rect 459560 3340 459612 3392
rect 460848 3340 460900 3392
rect 281264 3272 281316 3324
rect 288164 3272 288216 3324
rect 328828 3272 328880 3324
rect 333888 3272 333940 3324
rect 443000 3272 443052 3324
rect 232504 3204 232556 3256
rect 224132 3136 224184 3188
rect 232412 3136 232464 3188
rect 236000 3204 236052 3256
rect 251456 3204 251508 3256
rect 254584 3204 254636 3256
rect 253848 3136 253900 3188
rect 257068 3136 257120 3188
rect 243544 3068 243596 3120
rect 250352 3068 250404 3120
rect 251088 3068 251140 3120
rect 268936 3068 268988 3120
rect 280068 3204 280120 3256
rect 285588 3204 285640 3256
rect 286968 3136 287020 3188
rect 321652 3204 321704 3256
rect 322848 3204 322900 3256
rect 331128 3204 331180 3256
rect 435824 3204 435876 3256
rect 324044 3136 324096 3188
rect 328368 3136 328420 3188
rect 428740 3136 428792 3188
rect 285496 3068 285548 3120
rect 321652 3068 321704 3120
rect 262864 3000 262916 3052
rect 264612 3000 264664 3052
rect 284116 3000 284168 3052
rect 320456 3000 320508 3052
rect 325608 3068 325660 3120
rect 322756 3000 322808 3052
rect 414480 3000 414532 3052
rect 416780 3068 416832 3120
rect 417976 3068 418028 3120
rect 421564 3000 421616 3052
rect 10048 2932 10100 2984
rect 11704 2932 11756 2984
rect 24308 2932 24360 2984
rect 28264 2932 28316 2984
rect 113548 2932 113600 2984
rect 114468 2932 114520 2984
rect 120632 2932 120684 2984
rect 121368 2932 121420 2984
rect 114744 2864 114796 2916
rect 103980 2796 104032 2848
rect 107568 2796 107620 2848
rect 197636 2932 197688 2984
rect 231308 2932 231360 2984
rect 235264 2932 235316 2984
rect 263508 2932 263560 2984
rect 269304 2932 269356 2984
rect 282736 2932 282788 2984
rect 316960 2932 317012 2984
rect 317328 2932 317380 2984
rect 200304 2864 200356 2916
rect 245568 2864 245620 2916
rect 246304 2864 246356 2916
rect 284208 2864 284260 2916
rect 318064 2864 318116 2916
rect 325240 2932 325292 2984
rect 320088 2864 320140 2916
rect 407304 2932 407356 2984
rect 400220 2864 400272 2916
rect 121828 2796 121880 2848
rect 122748 2796 122800 2848
rect 124220 2796 124272 2848
rect 125508 2796 125560 2848
rect 125416 2728 125468 2780
rect 127808 2796 127860 2848
rect 128268 2796 128320 2848
rect 130200 2796 130252 2848
rect 131028 2796 131080 2848
rect 131396 2796 131448 2848
rect 132316 2796 132368 2848
rect 204260 2796 204312 2848
rect 255228 2796 255280 2848
rect 256240 2796 256292 2848
rect 256608 2796 256660 2848
rect 282828 2796 282880 2848
rect 314568 2796 314620 2848
rect 314660 2796 314712 2848
rect 393044 2796 393096 2848
rect 385132 2592 385184 2644
rect 385868 2592 385920 2644
rect 195612 1844 195664 1896
rect 205088 1232 205140 1284
rect 137284 552 137336 604
rect 137928 552 137980 604
rect 138480 552 138532 604
rect 139308 552 139360 604
rect 145656 552 145708 604
rect 146208 552 146260 604
rect 148048 552 148100 604
rect 148968 552 149020 604
rect 149244 552 149296 604
rect 150348 552 150400 604
rect 151544 552 151596 604
rect 151728 552 151780 604
rect 156328 552 156380 604
rect 157248 552 157300 604
rect 187240 552 187292 604
rect 187608 552 187660 604
rect 255044 595 255096 604
rect 255044 561 255053 595
rect 255053 561 255087 595
rect 255087 561 255096 595
rect 255044 552 255096 561
rect 259644 552 259696 604
rect 259828 552 259880 604
rect 265256 552 265308 604
rect 265808 552 265860 604
rect 300860 552 300912 604
rect 301412 552 301464 604
rect 307760 552 307812 604
rect 308588 552 308640 604
rect 309140 552 309192 604
rect 309784 552 309836 604
rect 314752 552 314804 604
rect 315764 552 315816 604
rect 325700 552 325752 604
rect 326436 552 326488 604
rect 332600 552 332652 604
rect 333612 552 333664 604
rect 336740 552 336792 604
rect 337108 552 337160 604
rect 339592 552 339644 604
rect 340696 552 340748 604
rect 378140 552 378192 604
rect 378784 552 378836 604
rect 520372 552 520424 604
rect 521476 552 521528 604
rect 524420 552 524472 604
rect 525064 552 525116 604
rect 531320 552 531372 604
rect 532240 552 532292 604
rect 538220 552 538272 604
rect 539324 552 539376 604
rect 542360 552 542412 604
rect 542912 552 542964 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 703474 8156 703520
rect 8036 703446 8156 703474
rect 8036 698290 8064 703446
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 72988 703474 73016 703520
rect 72804 703446 73016 703474
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 8024 698284 8076 698290
rect 8024 698226 8076 698232
rect 8208 698284 8260 698290
rect 8208 698226 8260 698232
rect 8220 695502 8248 698226
rect 8208 695496 8260 695502
rect 8208 695438 8260 695444
rect 8116 685908 8168 685914
rect 8116 685850 8168 685856
rect 3330 682272 3386 682281
rect 3330 682207 3386 682216
rect 3344 681766 3372 682207
rect 3332 681760 3384 681766
rect 3332 681702 3384 681708
rect 6184 681760 6236 681766
rect 6184 681702 6236 681708
rect 3422 667992 3478 668001
rect 3422 667927 3478 667936
rect 3054 624880 3110 624889
rect 3054 624815 3110 624824
rect 3068 623830 3096 624815
rect 3056 623824 3108 623830
rect 3056 623766 3108 623772
rect 3330 509960 3386 509969
rect 3330 509895 3386 509904
rect 3344 509794 3372 509895
rect 3332 509788 3384 509794
rect 3332 509730 3384 509736
rect 3330 452432 3386 452441
rect 3330 452367 3386 452376
rect 3344 451450 3372 452367
rect 3332 451444 3384 451450
rect 3332 451386 3384 451392
rect 3330 438016 3386 438025
rect 3330 437951 3386 437960
rect 3344 437714 3372 437951
rect 3332 437708 3384 437714
rect 3332 437650 3384 437656
rect 3330 423736 3386 423745
rect 3330 423671 3386 423680
rect 3344 342242 3372 423671
rect 3436 404326 3464 667927
rect 3514 653576 3570 653585
rect 3514 653511 3570 653520
rect 3528 409834 3556 653511
rect 3606 610464 3662 610473
rect 3606 610399 3662 610408
rect 3516 409828 3568 409834
rect 3516 409770 3568 409776
rect 3424 404320 3476 404326
rect 3424 404262 3476 404268
rect 3422 395040 3478 395049
rect 3422 394975 3478 394984
rect 3332 342236 3384 342242
rect 3332 342178 3384 342184
rect 3436 313274 3464 394975
rect 3620 386374 3648 610399
rect 3698 596048 3754 596057
rect 3698 595983 3754 595992
rect 3712 393310 3740 595983
rect 4066 567352 4122 567361
rect 4066 567287 4122 567296
rect 4080 567254 4108 567287
rect 4068 567248 4120 567254
rect 4068 567190 4120 567196
rect 3790 553072 3846 553081
rect 3790 553007 3846 553016
rect 3700 393304 3752 393310
rect 3700 393246 3752 393252
rect 3608 386368 3660 386374
rect 3608 386310 3660 386316
rect 3514 380624 3570 380633
rect 3514 380559 3570 380568
rect 3528 318782 3556 380559
rect 3804 369850 3832 553007
rect 3882 538656 3938 538665
rect 3882 538591 3938 538600
rect 3896 375358 3924 538591
rect 3974 495544 4030 495553
rect 3974 495479 4030 495488
rect 3884 375352 3936 375358
rect 3884 375294 3936 375300
rect 3792 369844 3844 369850
rect 3792 369786 3844 369792
rect 3606 366208 3662 366217
rect 3606 366143 3662 366152
rect 3620 324290 3648 366143
rect 3988 353258 4016 495479
rect 4066 481128 4122 481137
rect 4066 481063 4122 481072
rect 4080 358766 4108 481063
rect 4804 437708 4856 437714
rect 4804 437650 4856 437656
rect 4068 358760 4120 358766
rect 4068 358702 4120 358708
rect 3976 353252 4028 353258
rect 3976 353194 4028 353200
rect 3698 337512 3754 337521
rect 3698 337447 3754 337456
rect 3608 324284 3660 324290
rect 3608 324226 3660 324232
rect 3516 318776 3568 318782
rect 3516 318718 3568 318724
rect 3424 313268 3476 313274
rect 3424 313210 3476 313216
rect 3054 308816 3110 308825
rect 3054 308751 3110 308760
rect 3068 307766 3096 308751
rect 3056 307760 3108 307766
rect 3056 307702 3108 307708
rect 3712 296682 3740 337447
rect 4816 336734 4844 437650
rect 6196 398818 6224 681702
rect 8128 679046 8156 685850
rect 8116 679040 8168 679046
rect 8116 678982 8168 678988
rect 8024 678972 8076 678978
rect 8024 678914 8076 678920
rect 8036 673538 8064 678914
rect 8024 673532 8076 673538
rect 8024 673474 8076 673480
rect 8208 673532 8260 673538
rect 8208 673474 8260 673480
rect 8220 663762 8248 673474
rect 8036 663734 8248 663762
rect 8036 654158 8064 663734
rect 8024 654152 8076 654158
rect 8024 654094 8076 654100
rect 8208 654152 8260 654158
rect 8208 654094 8260 654100
rect 8220 644450 8248 654094
rect 8036 644422 8248 644450
rect 8036 634846 8064 644422
rect 8024 634840 8076 634846
rect 8024 634782 8076 634788
rect 8208 634840 8260 634846
rect 8208 634782 8260 634788
rect 8220 625138 8248 634782
rect 8036 625110 8248 625138
rect 8036 615534 8064 625110
rect 8024 615528 8076 615534
rect 8024 615470 8076 615476
rect 8208 615528 8260 615534
rect 8208 615470 8260 615476
rect 8220 605826 8248 615470
rect 8036 605798 8248 605826
rect 8036 596222 8064 605798
rect 8024 596216 8076 596222
rect 8208 596216 8260 596222
rect 8024 596158 8076 596164
rect 8128 596164 8208 596170
rect 8128 596158 8260 596164
rect 8128 596142 8248 596158
rect 8128 591954 8156 596142
rect 8036 591926 8156 591954
rect 8036 589286 8064 591926
rect 8024 589280 8076 589286
rect 8024 589222 8076 589228
rect 8024 579760 8076 579766
rect 7944 579708 8024 579714
rect 7944 579702 8076 579708
rect 7944 579686 8064 579702
rect 7944 579630 7972 579686
rect 7932 579624 7984 579630
rect 7932 579566 7984 579572
rect 8116 579624 8168 579630
rect 8116 579566 8168 579572
rect 8128 562970 8156 579566
rect 15844 567248 15896 567254
rect 15844 567190 15896 567196
rect 7932 562964 7984 562970
rect 7932 562906 7984 562912
rect 8116 562964 8168 562970
rect 8116 562906 8168 562912
rect 7944 553330 7972 562906
rect 7944 553302 8064 553330
rect 8036 550594 8064 553302
rect 8024 550588 8076 550594
rect 8024 550530 8076 550536
rect 8208 541000 8260 541006
rect 8208 540942 8260 540948
rect 8220 534018 8248 540942
rect 8128 533990 8248 534018
rect 8128 531321 8156 533990
rect 8114 531312 8170 531321
rect 8114 531247 8170 531256
rect 8390 531312 8446 531321
rect 8390 531247 8446 531256
rect 8404 521694 8432 531247
rect 8208 521688 8260 521694
rect 8208 521630 8260 521636
rect 8392 521688 8444 521694
rect 8392 521630 8444 521636
rect 8220 514706 8248 521630
rect 8128 514678 8248 514706
rect 8128 512009 8156 514678
rect 8114 512000 8170 512009
rect 8114 511935 8170 511944
rect 8390 512000 8446 512009
rect 8390 511935 8446 511944
rect 8404 502382 8432 511935
rect 10324 509788 10376 509794
rect 10324 509730 10376 509736
rect 8208 502376 8260 502382
rect 8208 502318 8260 502324
rect 8392 502376 8444 502382
rect 8392 502318 8444 502324
rect 8220 495394 8248 502318
rect 8128 495366 8248 495394
rect 8128 485858 8156 495366
rect 8116 485852 8168 485858
rect 8116 485794 8168 485800
rect 8208 485784 8260 485790
rect 8208 485726 8260 485732
rect 8220 483002 8248 485726
rect 7932 482996 7984 483002
rect 7932 482938 7984 482944
rect 8208 482996 8260 483002
rect 8208 482938 8260 482944
rect 7944 473385 7972 482938
rect 7930 473376 7986 473385
rect 7930 473311 7986 473320
rect 8114 473376 8170 473385
rect 8114 473311 8170 473320
rect 8128 466478 8156 473311
rect 8116 466472 8168 466478
rect 8116 466414 8168 466420
rect 8208 466404 8260 466410
rect 8208 466346 8260 466352
rect 8220 456770 8248 466346
rect 8036 456742 8248 456770
rect 8036 454034 8064 456742
rect 8024 454028 8076 454034
rect 8024 453970 8076 453976
rect 7932 444440 7984 444446
rect 7932 444382 7984 444388
rect 7944 437458 7972 444382
rect 7944 437430 8064 437458
rect 8036 427854 8064 437430
rect 8024 427848 8076 427854
rect 8024 427790 8076 427796
rect 8116 427780 8168 427786
rect 8116 427722 8168 427728
rect 8128 425066 8156 427722
rect 7840 425060 7892 425066
rect 7840 425002 7892 425008
rect 8116 425060 8168 425066
rect 8116 425002 8168 425008
rect 7852 415449 7880 425002
rect 7838 415440 7894 415449
rect 7838 415375 7894 415384
rect 8022 415440 8078 415449
rect 8022 415375 8078 415384
rect 8036 414730 8064 415375
rect 8024 414724 8076 414730
rect 8024 414666 8076 414672
rect 6184 398812 6236 398818
rect 6184 398754 6236 398760
rect 10336 347750 10364 509730
rect 11704 451444 11756 451450
rect 11704 451386 11756 451392
rect 10324 347744 10376 347750
rect 10324 347686 10376 347692
rect 4804 336728 4856 336734
rect 4804 336670 4856 336676
rect 11716 331226 11744 451386
rect 15856 364342 15884 567190
rect 24780 414798 24808 699654
rect 41340 414866 41368 700334
rect 72804 698306 72832 703446
rect 89180 699718 89208 703520
rect 105464 699718 105492 703520
rect 137848 703474 137876 703520
rect 137756 703446 137876 703474
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 89628 699712 89680 699718
rect 89628 699654 89680 699660
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 72712 698278 72832 698306
rect 72712 694142 72740 698278
rect 72700 694136 72752 694142
rect 72700 694078 72752 694084
rect 72516 684616 72568 684622
rect 72516 684558 72568 684564
rect 72528 684486 72556 684558
rect 72516 684480 72568 684486
rect 72516 684422 72568 684428
rect 72792 676116 72844 676122
rect 72792 676058 72844 676064
rect 72804 669390 72832 676058
rect 72792 669384 72844 669390
rect 72792 669326 72844 669332
rect 72792 669248 72844 669254
rect 72792 669190 72844 669196
rect 72804 659682 72832 669190
rect 72804 659666 72924 659682
rect 72804 659660 72936 659666
rect 72804 659654 72884 659660
rect 72884 659602 72936 659608
rect 73068 659660 73120 659666
rect 73068 659602 73120 659608
rect 73080 656878 73108 659602
rect 73068 656872 73120 656878
rect 73068 656814 73120 656820
rect 72976 647284 73028 647290
rect 72976 647226 73028 647232
rect 72988 640422 73016 647226
rect 72976 640416 73028 640422
rect 72976 640358 73028 640364
rect 72792 640280 72844 640286
rect 72792 640222 72844 640228
rect 72804 637566 72832 640222
rect 72792 637560 72844 637566
rect 72792 637502 72844 637508
rect 72884 637560 72936 637566
rect 72884 637502 72936 637508
rect 72896 630578 72924 637502
rect 72896 630550 73108 630578
rect 73080 626550 73108 630550
rect 73068 626544 73120 626550
rect 73068 626486 73120 626492
rect 73068 616888 73120 616894
rect 73068 616830 73120 616836
rect 73080 611454 73108 616830
rect 73068 611448 73120 611454
rect 73068 611390 73120 611396
rect 72884 611312 72936 611318
rect 72884 611254 72936 611260
rect 72896 608546 72924 611254
rect 72974 608560 73030 608569
rect 72896 608518 72974 608546
rect 72974 608495 73030 608504
rect 73158 608560 73214 608569
rect 73158 608495 73214 608504
rect 73172 601594 73200 608495
rect 72976 601588 73028 601594
rect 72976 601530 73028 601536
rect 73160 601588 73212 601594
rect 73160 601530 73212 601536
rect 72988 598942 73016 601530
rect 72976 598936 73028 598942
rect 72976 598878 73028 598884
rect 72884 589348 72936 589354
rect 72884 589290 72936 589296
rect 72896 582418 72924 589290
rect 72700 582412 72752 582418
rect 72700 582354 72752 582360
rect 72884 582412 72936 582418
rect 72884 582354 72936 582360
rect 72712 579630 72740 582354
rect 72700 579624 72752 579630
rect 72700 579566 72752 579572
rect 72608 569968 72660 569974
rect 72608 569910 72660 569916
rect 72620 563106 72648 569910
rect 72608 563100 72660 563106
rect 72608 563042 72660 563048
rect 72700 562964 72752 562970
rect 72700 562906 72752 562912
rect 72712 560266 72740 562906
rect 72620 560238 72740 560266
rect 72620 553450 72648 560238
rect 72608 553444 72660 553450
rect 72608 553386 72660 553392
rect 72608 550656 72660 550662
rect 72608 550598 72660 550604
rect 72620 543794 72648 550598
rect 72608 543788 72660 543794
rect 72608 543730 72660 543736
rect 72700 543652 72752 543658
rect 72700 543594 72752 543600
rect 72712 540954 72740 543594
rect 72620 540926 72740 540954
rect 72620 534138 72648 540926
rect 72608 534132 72660 534138
rect 72608 534074 72660 534080
rect 72620 531350 72648 531381
rect 72608 531344 72660 531350
rect 72698 531312 72754 531321
rect 72660 531292 72698 531298
rect 72608 531286 72698 531292
rect 72620 531270 72698 531286
rect 72698 531247 72754 531256
rect 72882 531312 72938 531321
rect 72882 531247 72938 531256
rect 72896 524346 72924 531247
rect 72700 524340 72752 524346
rect 72700 524282 72752 524288
rect 72884 524340 72936 524346
rect 72884 524282 72936 524288
rect 72712 514706 72740 524282
rect 72712 514678 72832 514706
rect 72804 512009 72832 514678
rect 72606 512000 72662 512009
rect 72606 511935 72662 511944
rect 72790 512000 72846 512009
rect 72790 511935 72846 511944
rect 72620 502382 72648 511935
rect 72608 502376 72660 502382
rect 72608 502318 72660 502324
rect 73068 502376 73120 502382
rect 73068 502318 73120 502324
rect 73080 495394 73108 502318
rect 72988 495366 73108 495394
rect 72988 485874 73016 495366
rect 72896 485846 73016 485874
rect 72896 480282 72924 485846
rect 72884 480276 72936 480282
rect 72884 480218 72936 480224
rect 73068 480276 73120 480282
rect 73068 480218 73120 480224
rect 73080 480162 73108 480218
rect 72988 480134 73108 480162
rect 72988 470642 73016 480134
rect 72896 470614 73016 470642
rect 72896 460970 72924 470614
rect 72884 460964 72936 460970
rect 72884 460906 72936 460912
rect 73068 460964 73120 460970
rect 73068 460906 73120 460912
rect 73080 460850 73108 460906
rect 72988 460822 73108 460850
rect 72988 444378 73016 460822
rect 72976 444372 73028 444378
rect 72976 444314 73028 444320
rect 73160 444372 73212 444378
rect 73160 444314 73212 444320
rect 73172 434761 73200 444314
rect 72882 434752 72938 434761
rect 72882 434687 72938 434696
rect 73158 434752 73214 434761
rect 73158 434687 73214 434696
rect 72896 425241 72924 434687
rect 72882 425232 72938 425241
rect 72882 425167 72938 425176
rect 72606 425096 72662 425105
rect 72662 425054 72740 425082
rect 72606 425031 72662 425040
rect 72712 418266 72740 425054
rect 72700 418260 72752 418266
rect 72700 418202 72752 418208
rect 72608 418124 72660 418130
rect 72608 418066 72660 418072
rect 72620 414934 72648 418066
rect 89640 415002 89668 699654
rect 106200 415070 106228 699654
rect 137756 698290 137784 703446
rect 137744 698284 137796 698290
rect 137744 698226 137796 698232
rect 137928 698284 137980 698290
rect 137928 698226 137980 698232
rect 137940 695502 137968 698226
rect 154132 695570 154160 703520
rect 170324 700262 170352 703520
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 171048 700256 171100 700262
rect 171048 700198 171100 700204
rect 154120 695564 154172 695570
rect 154120 695506 154172 695512
rect 154212 695564 154264 695570
rect 154212 695506 154264 695512
rect 137928 695496 137980 695502
rect 137928 695438 137980 695444
rect 154224 688634 154252 695506
rect 154212 688628 154264 688634
rect 154212 688570 154264 688576
rect 154396 688628 154448 688634
rect 154396 688570 154448 688576
rect 137836 685908 137888 685914
rect 137836 685850 137888 685856
rect 137848 679046 137876 685850
rect 154408 685846 154436 688570
rect 154396 685840 154448 685846
rect 154396 685782 154448 685788
rect 137836 679040 137888 679046
rect 137836 678982 137888 678988
rect 137744 678972 137796 678978
rect 137744 678914 137796 678920
rect 137756 673538 137784 678914
rect 154304 676252 154356 676258
rect 154304 676194 154356 676200
rect 154316 673538 154344 676194
rect 137744 673532 137796 673538
rect 137744 673474 137796 673480
rect 137928 673532 137980 673538
rect 137928 673474 137980 673480
rect 154304 673532 154356 673538
rect 154304 673474 154356 673480
rect 154488 673532 154540 673538
rect 154488 673474 154540 673480
rect 137940 663762 137968 673474
rect 154500 663762 154528 673474
rect 137756 663734 137968 663762
rect 154316 663734 154528 663762
rect 137756 654158 137784 663734
rect 154316 654158 154344 663734
rect 137744 654152 137796 654158
rect 137744 654094 137796 654100
rect 137928 654152 137980 654158
rect 137928 654094 137980 654100
rect 154304 654152 154356 654158
rect 154304 654094 154356 654100
rect 154488 654152 154540 654158
rect 154488 654094 154540 654100
rect 137940 644450 137968 654094
rect 154500 644450 154528 654094
rect 137756 644422 137968 644450
rect 154316 644422 154528 644450
rect 137756 634846 137784 644422
rect 154316 634846 154344 644422
rect 137744 634840 137796 634846
rect 137744 634782 137796 634788
rect 137928 634840 137980 634846
rect 137928 634782 137980 634788
rect 154304 634840 154356 634846
rect 154304 634782 154356 634788
rect 154488 634840 154540 634846
rect 154488 634782 154540 634788
rect 137940 625138 137968 634782
rect 154500 625138 154528 634782
rect 137756 625110 137968 625138
rect 154316 625110 154528 625138
rect 133144 623824 133196 623830
rect 133144 623766 133196 623772
rect 106188 415064 106240 415070
rect 106188 415006 106240 415012
rect 89628 414996 89680 415002
rect 89628 414938 89680 414944
rect 72608 414928 72660 414934
rect 72608 414870 72660 414876
rect 41328 414860 41380 414866
rect 41328 414802 41380 414808
rect 24768 414792 24820 414798
rect 24768 414734 24820 414740
rect 133156 380866 133184 623766
rect 137756 615534 137784 625110
rect 154316 615534 154344 625110
rect 137744 615528 137796 615534
rect 137744 615470 137796 615476
rect 137928 615528 137980 615534
rect 137928 615470 137980 615476
rect 154304 615528 154356 615534
rect 154304 615470 154356 615476
rect 154488 615528 154540 615534
rect 154488 615470 154540 615476
rect 137940 605826 137968 615470
rect 154500 605826 154528 615470
rect 137756 605798 137968 605826
rect 154316 605798 154528 605826
rect 137756 596222 137784 605798
rect 154316 596222 154344 605798
rect 137744 596216 137796 596222
rect 137928 596216 137980 596222
rect 137744 596158 137796 596164
rect 137848 596164 137928 596170
rect 137848 596158 137980 596164
rect 154304 596216 154356 596222
rect 154488 596216 154540 596222
rect 154304 596158 154356 596164
rect 154408 596164 154488 596170
rect 154408 596158 154540 596164
rect 137848 596142 137968 596158
rect 154408 596142 154528 596158
rect 137848 591954 137876 596142
rect 154408 591954 154436 596142
rect 137756 591926 137876 591954
rect 154316 591926 154436 591954
rect 137756 589286 137784 591926
rect 154316 589286 154344 591926
rect 137744 589280 137796 589286
rect 137744 589222 137796 589228
rect 154304 589280 154356 589286
rect 154304 589222 154356 589228
rect 137744 579760 137796 579766
rect 137664 579708 137744 579714
rect 154304 579760 154356 579766
rect 137664 579702 137796 579708
rect 154224 579708 154304 579714
rect 154224 579702 154356 579708
rect 137664 579686 137784 579702
rect 154224 579686 154344 579702
rect 137664 579630 137692 579686
rect 154224 579630 154252 579686
rect 137652 579624 137704 579630
rect 137652 579566 137704 579572
rect 154212 579624 154264 579630
rect 154212 579566 154264 579572
rect 154396 579624 154448 579630
rect 154396 579566 154448 579572
rect 137560 569968 137612 569974
rect 137560 569910 137612 569916
rect 137572 563106 137600 569910
rect 137560 563100 137612 563106
rect 137560 563042 137612 563048
rect 154408 562970 154436 579566
rect 137652 562964 137704 562970
rect 137652 562906 137704 562912
rect 154212 562964 154264 562970
rect 154212 562906 154264 562912
rect 154396 562964 154448 562970
rect 154396 562906 154448 562912
rect 137664 560250 137692 562906
rect 137652 560244 137704 560250
rect 137652 560186 137704 560192
rect 154224 553330 154252 562906
rect 154224 553302 154344 553330
rect 137836 550656 137888 550662
rect 137836 550598 137888 550604
rect 137848 543658 137876 550598
rect 154316 543810 154344 553302
rect 154316 543782 154528 543810
rect 137652 543652 137704 543658
rect 137652 543594 137704 543600
rect 137836 543652 137888 543658
rect 137836 543594 137888 543600
rect 137664 534070 137692 543594
rect 137652 534064 137704 534070
rect 137652 534006 137704 534012
rect 137836 534064 137888 534070
rect 154500 534018 154528 543782
rect 137836 534006 137888 534012
rect 137848 531321 137876 534006
rect 154408 533990 154528 534018
rect 137834 531312 137890 531321
rect 137834 531247 137890 531256
rect 138110 531312 138166 531321
rect 154408 531282 154436 533990
rect 138110 531247 138166 531256
rect 154396 531276 154448 531282
rect 138124 521694 138152 531247
rect 154396 531218 154448 531224
rect 137928 521688 137980 521694
rect 137928 521630 137980 521636
rect 138112 521688 138164 521694
rect 138112 521630 138164 521636
rect 154488 521688 154540 521694
rect 154488 521630 154540 521636
rect 137940 514706 137968 521630
rect 154500 514706 154528 521630
rect 137848 514678 137968 514706
rect 154408 514678 154528 514706
rect 137848 512009 137876 514678
rect 137834 512000 137890 512009
rect 137834 511935 137890 511944
rect 138110 512000 138166 512009
rect 154408 511970 154436 514678
rect 138110 511935 138166 511944
rect 154396 511964 154448 511970
rect 138124 502382 138152 511935
rect 154396 511906 154448 511912
rect 137928 502376 137980 502382
rect 137928 502318 137980 502324
rect 138112 502376 138164 502382
rect 138112 502318 138164 502324
rect 154488 502376 154540 502382
rect 154488 502318 154540 502324
rect 137940 495394 137968 502318
rect 154500 495394 154528 502318
rect 137848 495366 137968 495394
rect 154408 495366 154528 495394
rect 137848 492658 137876 495366
rect 154408 492658 154436 495366
rect 137652 492652 137704 492658
rect 137652 492594 137704 492600
rect 137836 492652 137888 492658
rect 137836 492594 137888 492600
rect 154212 492652 154264 492658
rect 154212 492594 154264 492600
rect 154396 492652 154448 492658
rect 154396 492594 154448 492600
rect 137664 483041 137692 492594
rect 154224 483041 154252 492594
rect 137650 483032 137706 483041
rect 137650 482967 137706 482976
rect 137926 483032 137982 483041
rect 137926 482967 137982 482976
rect 154210 483032 154266 483041
rect 154210 482967 154266 482976
rect 154486 483032 154542 483041
rect 154486 482967 154542 482976
rect 137940 476082 137968 482967
rect 154500 476082 154528 482967
rect 137756 476054 137968 476082
rect 154316 476054 154528 476082
rect 137756 466546 137784 476054
rect 137744 466540 137796 466546
rect 137744 466482 137796 466488
rect 154316 466478 154344 476054
rect 154304 466472 154356 466478
rect 154304 466414 154356 466420
rect 154488 466472 154540 466478
rect 154488 466414 154540 466420
rect 137652 466404 137704 466410
rect 137652 466346 137704 466352
rect 137664 463690 137692 466346
rect 137376 463684 137428 463690
rect 137376 463626 137428 463632
rect 137652 463684 137704 463690
rect 137652 463626 137704 463632
rect 137388 454073 137416 463626
rect 154500 456770 154528 466414
rect 154316 456742 154528 456770
rect 137374 454064 137430 454073
rect 137374 453999 137430 454008
rect 137558 454064 137614 454073
rect 154316 454034 154344 456742
rect 137558 453999 137614 454008
rect 154304 454028 154356 454034
rect 137572 447166 137600 453999
rect 154304 453970 154356 453976
rect 137560 447160 137612 447166
rect 137560 447102 137612 447108
rect 137652 447092 137704 447098
rect 137652 447034 137704 447040
rect 137664 437458 137692 447034
rect 154212 444440 154264 444446
rect 154212 444382 154264 444388
rect 154224 437458 154252 444382
rect 137664 437430 137784 437458
rect 154224 437430 154344 437458
rect 137756 427854 137784 437430
rect 154316 427854 154344 437430
rect 137744 427848 137796 427854
rect 137744 427790 137796 427796
rect 154304 427848 154356 427854
rect 154304 427790 154356 427796
rect 137836 427780 137888 427786
rect 137836 427722 137888 427728
rect 154396 427780 154448 427786
rect 154396 427722 154448 427728
rect 137848 425066 137876 427722
rect 154408 425066 154436 427722
rect 137560 425060 137612 425066
rect 137560 425002 137612 425008
rect 137836 425060 137888 425066
rect 137836 425002 137888 425008
rect 154120 425060 154172 425066
rect 154120 425002 154172 425008
rect 154396 425060 154448 425066
rect 154396 425002 154448 425008
rect 137572 415449 137600 425002
rect 154132 415449 154160 425002
rect 137558 415440 137614 415449
rect 137558 415375 137614 415384
rect 137742 415440 137798 415449
rect 137742 415375 137798 415384
rect 154118 415440 154174 415449
rect 154118 415375 154174 415384
rect 154302 415440 154358 415449
rect 154302 415375 154358 415384
rect 137756 415138 137784 415375
rect 154316 415206 154344 415375
rect 154304 415200 154356 415206
rect 154304 415142 154356 415148
rect 137744 415132 137796 415138
rect 137744 415074 137796 415080
rect 168012 414792 168064 414798
rect 168012 414734 168064 414740
rect 159364 414724 159416 414730
rect 159364 414666 159416 414672
rect 159376 411740 159404 414666
rect 168024 411740 168052 414734
rect 171060 414730 171088 700198
rect 202420 415064 202472 415070
rect 202420 415006 202472 415012
rect 194048 414996 194100 415002
rect 194048 414938 194100 414944
rect 185400 414928 185452 414934
rect 185400 414870 185452 414876
rect 176660 414860 176712 414866
rect 176660 414802 176712 414808
rect 171048 414724 171100 414730
rect 171048 414666 171100 414672
rect 176672 411740 176700 414802
rect 185412 411740 185440 414870
rect 194060 411740 194088 414938
rect 202432 411754 202460 415006
rect 202800 414798 202828 703520
rect 218992 703474 219020 703520
rect 218900 703446 219020 703474
rect 218900 695745 218928 703446
rect 235184 699718 235212 703520
rect 267660 699718 267688 703520
rect 283852 700398 283880 703520
rect 289728 700460 289780 700466
rect 289728 700402 289780 700408
rect 273168 700392 273220 700398
rect 273168 700334 273220 700340
rect 283840 700392 283892 700398
rect 283840 700334 283892 700340
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 264888 699712 264940 699718
rect 264888 699654 264940 699660
rect 267648 699712 267700 699718
rect 267648 699654 267700 699660
rect 218886 695736 218942 695745
rect 218886 695671 218942 695680
rect 219254 695600 219310 695609
rect 219176 695558 219254 695586
rect 219176 695502 219204 695558
rect 219254 695535 219310 695544
rect 219164 695496 219216 695502
rect 219164 695438 219216 695444
rect 219072 685908 219124 685914
rect 219072 685850 219124 685856
rect 219084 678994 219112 685850
rect 218992 678966 219112 678994
rect 218992 676190 219020 678966
rect 218980 676184 219032 676190
rect 218980 676126 219032 676132
rect 219072 666596 219124 666602
rect 219072 666538 219124 666544
rect 219084 659682 219112 666538
rect 219084 659666 219204 659682
rect 219084 659660 219216 659666
rect 219084 659654 219164 659660
rect 219164 659602 219216 659608
rect 219348 659660 219400 659666
rect 219348 659602 219400 659608
rect 219360 656878 219388 659602
rect 219348 656872 219400 656878
rect 219348 656814 219400 656820
rect 219256 647284 219308 647290
rect 219256 647226 219308 647232
rect 219268 640422 219296 647226
rect 219256 640416 219308 640422
rect 219256 640358 219308 640364
rect 219072 640280 219124 640286
rect 219072 640222 219124 640228
rect 219084 637566 219112 640222
rect 219072 637560 219124 637566
rect 219072 637502 219124 637508
rect 219164 637560 219216 637566
rect 219164 637502 219216 637508
rect 219176 630578 219204 637502
rect 219176 630550 219388 630578
rect 219360 626550 219388 630550
rect 219348 626544 219400 626550
rect 219348 626486 219400 626492
rect 219348 616888 219400 616894
rect 219348 616830 219400 616836
rect 219360 611454 219388 616830
rect 219348 611448 219400 611454
rect 219348 611390 219400 611396
rect 219072 608728 219124 608734
rect 219072 608670 219124 608676
rect 219084 608598 219112 608670
rect 219072 608592 219124 608598
rect 219072 608534 219124 608540
rect 219256 601588 219308 601594
rect 219256 601530 219308 601536
rect 219268 598942 219296 601530
rect 219256 598936 219308 598942
rect 219256 598878 219308 598884
rect 219164 589348 219216 589354
rect 219164 589290 219216 589296
rect 219176 582418 219204 589290
rect 218980 582412 219032 582418
rect 218980 582354 219032 582360
rect 219164 582412 219216 582418
rect 219164 582354 219216 582360
rect 218992 579630 219020 582354
rect 218980 579624 219032 579630
rect 218980 579566 219032 579572
rect 218888 569968 218940 569974
rect 218888 569910 218940 569916
rect 218900 563106 218928 569910
rect 218888 563100 218940 563106
rect 218888 563042 218940 563048
rect 218980 562964 219032 562970
rect 218980 562906 219032 562912
rect 218992 560266 219020 562906
rect 218900 560238 219020 560266
rect 218900 553450 218928 560238
rect 218888 553444 218940 553450
rect 218888 553386 218940 553392
rect 218888 550656 218940 550662
rect 218888 550598 218940 550604
rect 218900 543794 218928 550598
rect 218888 543788 218940 543794
rect 218888 543730 218940 543736
rect 218980 543652 219032 543658
rect 218980 543594 219032 543600
rect 218992 540977 219020 543594
rect 218978 540968 219034 540977
rect 218978 540903 219034 540912
rect 219162 540968 219218 540977
rect 219162 540903 219218 540912
rect 219176 533882 219204 540903
rect 218992 533854 219204 533882
rect 218992 531321 219020 533854
rect 218978 531312 219034 531321
rect 218978 531247 219034 531256
rect 219162 531312 219218 531321
rect 219162 531247 219218 531256
rect 219176 524346 219204 531247
rect 218980 524340 219032 524346
rect 218980 524282 219032 524288
rect 219164 524340 219216 524346
rect 219164 524282 219216 524288
rect 218992 514706 219020 524282
rect 218992 514678 219112 514706
rect 219084 512009 219112 514678
rect 218886 512000 218942 512009
rect 218886 511935 218942 511944
rect 219070 512000 219126 512009
rect 219070 511935 219126 511944
rect 218900 502382 218928 511935
rect 218888 502376 218940 502382
rect 218888 502318 218940 502324
rect 219348 502376 219400 502382
rect 219348 502318 219400 502324
rect 219360 495394 219388 502318
rect 219268 495366 219388 495394
rect 219268 485874 219296 495366
rect 219176 485846 219296 485874
rect 219176 480282 219204 485846
rect 219164 480276 219216 480282
rect 219164 480218 219216 480224
rect 219348 480276 219400 480282
rect 219348 480218 219400 480224
rect 219360 480162 219388 480218
rect 219268 480134 219388 480162
rect 219268 470642 219296 480134
rect 219176 470614 219296 470642
rect 219176 460970 219204 470614
rect 219164 460964 219216 460970
rect 219164 460906 219216 460912
rect 219348 460964 219400 460970
rect 219348 460906 219400 460912
rect 219360 460850 219388 460906
rect 219268 460822 219388 460850
rect 219268 444378 219296 460822
rect 219256 444372 219308 444378
rect 219256 444314 219308 444320
rect 219440 444372 219492 444378
rect 219440 444314 219492 444320
rect 219452 434761 219480 444314
rect 219162 434752 219218 434761
rect 219162 434687 219218 434696
rect 219438 434752 219494 434761
rect 219438 434687 219494 434696
rect 219176 425241 219204 434687
rect 219162 425232 219218 425241
rect 219162 425167 219218 425176
rect 218886 425096 218942 425105
rect 218942 425054 219020 425082
rect 218886 425031 218942 425040
rect 218992 418266 219020 425054
rect 218980 418260 219032 418266
rect 218980 418202 219032 418208
rect 218888 418124 218940 418130
rect 218888 418066 218940 418072
rect 211436 415132 211488 415138
rect 211436 415074 211488 415080
rect 202788 414792 202840 414798
rect 202788 414734 202840 414740
rect 202432 411726 202814 411754
rect 211448 411740 211476 415074
rect 218900 414866 218928 418066
rect 220176 415200 220228 415206
rect 220176 415142 220228 415148
rect 218888 414860 218940 414866
rect 218888 414802 218940 414808
rect 220188 411740 220216 415142
rect 235920 414730 235948 699654
rect 264900 415410 264928 699654
rect 263600 415404 263652 415410
rect 263600 415346 263652 415352
rect 264888 415404 264940 415410
rect 264888 415346 264940 415352
rect 246212 414860 246264 414866
rect 246212 414802 246264 414808
rect 237564 414792 237616 414798
rect 237564 414734 237616 414740
rect 228824 414724 228876 414730
rect 228824 414666 228876 414672
rect 235908 414724 235960 414730
rect 235908 414666 235960 414672
rect 228836 411740 228864 414666
rect 237576 411740 237604 414734
rect 246224 411740 246252 414802
rect 254952 414724 255004 414730
rect 254952 414666 255004 414672
rect 254964 411740 254992 414666
rect 263612 411740 263640 415346
rect 273180 414730 273208 700334
rect 281448 700324 281500 700330
rect 281448 700266 281500 700272
rect 272340 414724 272392 414730
rect 272340 414666 272392 414672
rect 273168 414724 273220 414730
rect 273168 414666 273220 414672
rect 272352 411740 272380 414666
rect 281460 411618 281488 700266
rect 289740 411740 289768 700402
rect 299388 700392 299440 700398
rect 299388 700334 299440 700340
rect 299400 415410 299428 700334
rect 300136 700330 300164 703520
rect 315948 700868 316000 700874
rect 315948 700810 316000 700816
rect 300124 700324 300176 700330
rect 300124 700266 300176 700272
rect 307668 700324 307720 700330
rect 307668 700266 307720 700272
rect 298376 415404 298428 415410
rect 298376 415346 298428 415352
rect 299388 415404 299440 415410
rect 299388 415346 299440 415352
rect 298388 411740 298416 415346
rect 307680 411618 307708 700266
rect 315960 411754 315988 700810
rect 325608 700800 325660 700806
rect 325608 700742 325660 700748
rect 325620 414254 325648 700742
rect 332520 700466 332548 703520
rect 333888 700732 333940 700738
rect 333888 700674 333940 700680
rect 332508 700460 332560 700466
rect 332508 700402 332560 700408
rect 324504 414248 324556 414254
rect 324504 414190 324556 414196
rect 325608 414248 325660 414254
rect 325608 414190 325660 414196
rect 315790 411726 315988 411754
rect 324516 411740 324544 414190
rect 333900 411618 333928 700674
rect 342168 700664 342220 700670
rect 342168 700606 342220 700612
rect 342180 411754 342208 700606
rect 348804 700398 348832 703520
rect 351828 700596 351880 700602
rect 351828 700538 351880 700544
rect 348792 700392 348844 700398
rect 348792 700334 348844 700340
rect 351840 415138 351868 700538
rect 360108 700528 360160 700534
rect 360108 700470 360160 700476
rect 360120 415410 360148 700470
rect 364996 700330 365024 703520
rect 397472 700874 397500 703520
rect 397460 700868 397512 700874
rect 397460 700810 397512 700816
rect 413664 700806 413692 703520
rect 413652 700800 413704 700806
rect 413652 700742 413704 700748
rect 429856 700738 429884 703520
rect 429844 700732 429896 700738
rect 429844 700674 429896 700680
rect 462332 700670 462360 703520
rect 462320 700664 462372 700670
rect 462320 700606 462372 700612
rect 478524 700602 478552 703520
rect 478512 700596 478564 700602
rect 478512 700538 478564 700544
rect 494808 700534 494836 703520
rect 494796 700528 494848 700534
rect 494796 700470 494848 700476
rect 527192 700466 527220 703520
rect 368388 700460 368440 700466
rect 368388 700402 368440 700408
rect 527180 700460 527232 700466
rect 527180 700402 527232 700408
rect 364984 700324 365036 700330
rect 364984 700266 365036 700272
rect 359280 415404 359332 415410
rect 359280 415346 359332 415352
rect 360108 415404 360160 415410
rect 360108 415346 360160 415352
rect 350540 415132 350592 415138
rect 350540 415074 350592 415080
rect 351828 415132 351880 415138
rect 351828 415074 351880 415080
rect 341918 411726 342208 411754
rect 350552 411740 350580 415074
rect 359292 411740 359320 415346
rect 368400 411754 368428 700402
rect 543476 700398 543504 703520
rect 376668 700392 376720 700398
rect 376668 700334 376720 700340
rect 543464 700392 543516 700398
rect 543464 700334 543516 700340
rect 367954 411726 368428 411754
rect 376680 411740 376708 700334
rect 559668 700330 559696 703520
rect 386328 700324 386380 700330
rect 386328 700266 386380 700272
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 386340 415410 386368 700266
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 393964 696992 394016 696998
rect 393964 696934 394016 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 392584 685908 392636 685914
rect 392584 685850 392636 685856
rect 385316 415404 385368 415410
rect 385316 415346 385368 415352
rect 386328 415404 386380 415410
rect 386328 415346 386380 415352
rect 385328 411740 385356 415346
rect 281014 411590 281488 411618
rect 307142 411590 307708 411618
rect 333178 411590 333928 411618
rect 151820 409828 151872 409834
rect 151820 409770 151872 409776
rect 151832 408921 151860 409770
rect 391940 409284 391992 409290
rect 391940 409226 391992 409232
rect 391952 409193 391980 409226
rect 391938 409184 391994 409193
rect 391938 409119 391994 409128
rect 151818 408912 151874 408921
rect 151818 408847 151874 408856
rect 152372 404320 152424 404326
rect 152372 404262 152424 404268
rect 152384 403345 152412 404262
rect 392596 403889 392624 685850
rect 392676 592068 392728 592074
rect 392676 592010 392728 592016
rect 392582 403880 392638 403889
rect 392582 403815 392638 403824
rect 152370 403336 152426 403345
rect 152370 403271 152426 403280
rect 153108 398812 153160 398818
rect 153108 398754 153160 398760
rect 391940 398812 391992 398818
rect 391940 398754 391992 398760
rect 153120 397633 153148 398754
rect 391952 398585 391980 398754
rect 391938 398576 391994 398585
rect 391938 398511 391994 398520
rect 153106 397624 153162 397633
rect 153106 397559 153162 397568
rect 391940 394664 391992 394670
rect 391940 394606 391992 394612
rect 391952 393417 391980 394606
rect 391938 393408 391994 393417
rect 391938 393343 391994 393352
rect 153108 393304 153160 393310
rect 153108 393246 153160 393252
rect 153120 392057 153148 393246
rect 153106 392048 153162 392057
rect 153106 391983 153162 391992
rect 391940 389156 391992 389162
rect 391940 389098 391992 389104
rect 391952 388113 391980 389098
rect 391938 388104 391994 388113
rect 391938 388039 391994 388048
rect 153108 386368 153160 386374
rect 153106 386336 153108 386345
rect 153160 386336 153162 386345
rect 153106 386271 153162 386280
rect 391940 383648 391992 383654
rect 391940 383590 391992 383596
rect 391952 382809 391980 383590
rect 391938 382800 391994 382809
rect 391938 382735 391994 382744
rect 133144 380860 133196 380866
rect 133144 380802 133196 380808
rect 152556 380860 152608 380866
rect 152556 380802 152608 380808
rect 152568 380769 152596 380802
rect 152554 380760 152610 380769
rect 152554 380695 152610 380704
rect 391940 378140 391992 378146
rect 391940 378082 391992 378088
rect 391952 377641 391980 378082
rect 391938 377632 391994 377641
rect 391938 377567 391994 377576
rect 152556 375352 152608 375358
rect 152556 375294 152608 375300
rect 152568 375057 152596 375294
rect 152554 375048 152610 375057
rect 152554 374983 152610 374992
rect 392688 372337 392716 592010
rect 392768 498228 392820 498234
rect 392768 498170 392820 498176
rect 392674 372328 392730 372337
rect 392674 372263 392730 372272
rect 152924 369844 152976 369850
rect 152924 369786 152976 369792
rect 152936 369481 152964 369786
rect 152922 369472 152978 369481
rect 152922 369407 152978 369416
rect 392584 368552 392636 368558
rect 392584 368494 392636 368500
rect 391940 367056 391992 367062
rect 391938 367024 391940 367033
rect 391992 367024 391994 367033
rect 391938 366959 391994 366968
rect 15844 364336 15896 364342
rect 15844 364278 15896 364284
rect 153108 364336 153160 364342
rect 153108 364278 153160 364284
rect 153120 363769 153148 364278
rect 153106 363760 153162 363769
rect 153106 363695 153162 363704
rect 391940 362908 391992 362914
rect 391940 362850 391992 362856
rect 391952 361865 391980 362850
rect 391938 361856 391994 361865
rect 391938 361791 391994 361800
rect 153108 358760 153160 358766
rect 153108 358702 153160 358708
rect 153120 358193 153148 358702
rect 153106 358184 153162 358193
rect 153106 358119 153162 358128
rect 391940 357400 391992 357406
rect 391940 357342 391992 357348
rect 391952 356561 391980 357342
rect 391938 356552 391994 356561
rect 391938 356487 391994 356496
rect 153108 353252 153160 353258
rect 153108 353194 153160 353200
rect 153120 352617 153148 353194
rect 153106 352608 153162 352617
rect 153106 352543 153162 352552
rect 391940 351892 391992 351898
rect 391940 351834 391992 351840
rect 391952 351257 391980 351834
rect 391938 351248 391994 351257
rect 391938 351183 391994 351192
rect 152924 347744 152976 347750
rect 152924 347686 152976 347692
rect 152936 346905 152964 347686
rect 152922 346896 152978 346905
rect 152922 346831 152978 346840
rect 391940 346384 391992 346390
rect 391940 346326 391992 346332
rect 391952 346089 391980 346326
rect 391938 346080 391994 346089
rect 391938 346015 391994 346024
rect 152556 342236 152608 342242
rect 152556 342178 152608 342184
rect 152568 341329 152596 342178
rect 152554 341320 152610 341329
rect 152554 341255 152610 341264
rect 153108 336728 153160 336734
rect 153108 336670 153160 336676
rect 391940 336728 391992 336734
rect 391940 336670 391992 336676
rect 153120 335617 153148 336670
rect 153106 335608 153162 335617
rect 153106 335543 153162 335552
rect 391952 335481 391980 336670
rect 391938 335472 391994 335481
rect 391938 335407 391994 335416
rect 11704 331220 11756 331226
rect 11704 331162 11756 331168
rect 153108 331220 153160 331226
rect 153108 331162 153160 331168
rect 153120 330041 153148 331162
rect 391940 330404 391992 330410
rect 391940 330346 391992 330352
rect 391952 330177 391980 330346
rect 391938 330168 391994 330177
rect 391938 330103 391994 330112
rect 153106 330032 153162 330041
rect 153106 329967 153162 329976
rect 391940 325644 391992 325650
rect 391940 325586 391992 325592
rect 391952 325009 391980 325586
rect 391938 325000 391994 325009
rect 391938 324935 391994 324944
rect 153106 324320 153162 324329
rect 153106 324255 153108 324264
rect 153160 324255 153162 324264
rect 153108 324226 153160 324232
rect 3790 323096 3846 323105
rect 3790 323031 3846 323040
rect 3804 302190 3832 323031
rect 391940 320136 391992 320142
rect 391940 320078 391992 320084
rect 391952 319705 391980 320078
rect 391938 319696 391994 319705
rect 391938 319631 391994 319640
rect 153108 318776 153160 318782
rect 153106 318744 153108 318753
rect 153160 318744 153162 318753
rect 153106 318679 153162 318688
rect 152372 313268 152424 313274
rect 152372 313210 152424 313216
rect 152384 313041 152412 313210
rect 152370 313032 152426 313041
rect 152370 312967 152426 312976
rect 391940 309596 391992 309602
rect 391940 309538 391992 309544
rect 391952 309233 391980 309538
rect 391938 309224 391994 309233
rect 391938 309159 391994 309168
rect 152556 307760 152608 307766
rect 152556 307702 152608 307708
rect 152568 307465 152596 307702
rect 152554 307456 152610 307465
rect 152554 307391 152610 307400
rect 391940 304972 391992 304978
rect 391940 304914 391992 304920
rect 391952 303929 391980 304914
rect 391938 303920 391994 303929
rect 391938 303855 391994 303864
rect 3792 302184 3844 302190
rect 3792 302126 3844 302132
rect 153108 302184 153160 302190
rect 153108 302126 153160 302132
rect 153120 301753 153148 302126
rect 153106 301744 153162 301753
rect 153106 301679 153162 301688
rect 392596 298625 392624 368494
rect 392676 357468 392728 357474
rect 392676 357410 392728 357416
rect 392582 298616 392638 298625
rect 392582 298551 392638 298560
rect 3700 296676 3752 296682
rect 3700 296618 3752 296624
rect 152740 296676 152792 296682
rect 152740 296618 152792 296624
rect 152752 296177 152780 296618
rect 152738 296168 152794 296177
rect 152738 296103 152794 296112
rect 3514 294400 3570 294409
rect 3514 294335 3570 294344
rect 3424 289876 3476 289882
rect 3424 289818 3476 289824
rect 2964 284368 3016 284374
rect 2964 284310 3016 284316
rect 2976 280129 3004 284310
rect 2962 280120 3018 280129
rect 2962 280055 3018 280064
rect 3436 265713 3464 289818
rect 3528 280158 3556 294335
rect 392688 293457 392716 357410
rect 392780 340785 392808 498170
rect 392860 415472 392912 415478
rect 392860 415414 392912 415420
rect 392766 340776 392822 340785
rect 392766 340711 392822 340720
rect 392768 321632 392820 321638
rect 392768 321574 392820 321580
rect 392674 293448 392730 293457
rect 392674 293383 392730 293392
rect 152186 290592 152242 290601
rect 152186 290527 152242 290536
rect 152200 289882 152228 290527
rect 152188 289876 152240 289882
rect 152188 289818 152240 289824
rect 391940 288380 391992 288386
rect 391940 288322 391992 288328
rect 391952 288153 391980 288322
rect 391938 288144 391994 288153
rect 391938 288079 391994 288088
rect 152002 284880 152058 284889
rect 152002 284815 152058 284824
rect 152016 284374 152044 284815
rect 152004 284368 152056 284374
rect 152004 284310 152056 284316
rect 392780 282849 392808 321574
rect 392872 314401 392900 415414
rect 393976 409290 394004 696934
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 580172 685850 580224 685856
rect 580262 674656 580318 674665
rect 580262 674591 580318 674600
rect 579894 639432 579950 639441
rect 579894 639367 579950 639376
rect 579908 638994 579936 639367
rect 398104 638988 398156 638994
rect 398104 638930 398156 638936
rect 579896 638988 579948 638994
rect 579896 638930 579948 638936
rect 396724 545148 396776 545154
rect 396724 545090 396776 545096
rect 395344 462392 395396 462398
rect 395344 462334 395396 462340
rect 393964 409284 394016 409290
rect 393964 409226 394016 409232
rect 393964 404388 394016 404394
rect 393964 404330 394016 404336
rect 392858 314392 392914 314401
rect 392858 314327 392914 314336
rect 392860 310548 392912 310554
rect 392860 310490 392912 310496
rect 392766 282840 392822 282849
rect 392766 282775 392822 282784
rect 3516 280152 3568 280158
rect 3516 280094 3568 280100
rect 152924 280152 152976 280158
rect 152924 280094 152976 280100
rect 152936 279313 152964 280094
rect 152922 279304 152978 279313
rect 152922 279239 152978 279248
rect 392872 277681 392900 310490
rect 393976 309602 394004 404330
rect 395356 330410 395384 462334
rect 396736 357406 396764 545090
rect 398116 389162 398144 638930
rect 580170 592512 580226 592521
rect 580170 592447 580226 592456
rect 580184 592074 580212 592447
rect 580172 592068 580224 592074
rect 580172 592010 580224 592016
rect 580170 545592 580226 545601
rect 580170 545527 580226 545536
rect 580184 545154 580212 545527
rect 580172 545148 580224 545154
rect 580172 545090 580224 545096
rect 579986 498672 580042 498681
rect 579986 498607 580042 498616
rect 580000 498234 580028 498607
rect 579988 498228 580040 498234
rect 579988 498170 580040 498176
rect 579986 486840 580042 486849
rect 579986 486775 580042 486784
rect 580000 485858 580028 486775
rect 400864 485852 400916 485858
rect 400864 485794 400916 485800
rect 579988 485852 580040 485858
rect 579988 485794 580040 485800
rect 399484 451308 399536 451314
rect 399484 451250 399536 451256
rect 398104 389156 398156 389162
rect 398104 389098 398156 389104
rect 396724 357400 396776 357406
rect 396724 357342 396776 357348
rect 395344 330404 395396 330410
rect 395344 330346 395396 330352
rect 399496 325650 399524 451250
rect 400876 336734 400904 485794
rect 579986 463448 580042 463457
rect 579986 463383 580042 463392
rect 580000 462398 580028 463383
rect 579988 462392 580040 462398
rect 579988 462334 580040 462340
rect 579986 451752 580042 451761
rect 579986 451687 580042 451696
rect 580000 451314 580028 451687
rect 579988 451308 580040 451314
rect 579988 451250 580040 451256
rect 580170 439920 580226 439929
rect 580170 439855 580226 439864
rect 580078 416528 580134 416537
rect 580078 416463 580134 416472
rect 580092 415478 580120 416463
rect 580080 415472 580132 415478
rect 580080 415414 580132 415420
rect 579896 412616 579948 412622
rect 579896 412558 579948 412564
rect 579908 404138 579936 412558
rect 580078 404832 580134 404841
rect 580078 404767 580134 404776
rect 580092 404394 580120 404767
rect 580080 404388 580132 404394
rect 580080 404330 580132 404336
rect 579908 404110 580120 404138
rect 580092 398818 580120 404110
rect 580080 398812 580132 398818
rect 580080 398754 580132 398760
rect 580078 369608 580134 369617
rect 580078 369543 580134 369552
rect 580092 368558 580120 369543
rect 580080 368552 580132 368558
rect 580080 368494 580132 368500
rect 580078 357912 580134 357921
rect 580078 357847 580134 357856
rect 580092 357474 580120 357847
rect 580080 357468 580132 357474
rect 580080 357410 580132 357416
rect 400864 336728 400916 336734
rect 400864 336670 400916 336676
rect 399484 325644 399536 325650
rect 399484 325586 399536 325592
rect 580184 322794 580212 439855
rect 580276 412622 580304 674591
rect 580354 651128 580410 651137
rect 580354 651063 580410 651072
rect 580264 412616 580316 412622
rect 580264 412558 580316 412564
rect 580368 394670 580396 651063
rect 580446 627736 580502 627745
rect 580446 627671 580502 627680
rect 580356 394664 580408 394670
rect 580356 394606 580408 394612
rect 580262 393000 580318 393009
rect 580262 392935 580318 392944
rect 579896 322788 579948 322794
rect 579896 322730 579948 322736
rect 580172 322788 580224 322794
rect 580172 322730 580224 322736
rect 579908 320142 579936 322730
rect 580170 322688 580226 322697
rect 580170 322623 580226 322632
rect 580184 321638 580212 322623
rect 580172 321632 580224 321638
rect 580172 321574 580224 321580
rect 579896 320136 579948 320142
rect 579896 320078 579948 320084
rect 579618 310856 579674 310865
rect 579618 310791 579674 310800
rect 579632 310554 579660 310791
rect 579620 310548 579672 310554
rect 579620 310490 579672 310496
rect 393964 309596 394016 309602
rect 393964 309538 394016 309544
rect 580276 304978 580304 392935
rect 580460 383654 580488 627671
rect 580538 604208 580594 604217
rect 580538 604143 580594 604152
rect 580448 383648 580500 383654
rect 580448 383590 580500 383596
rect 580552 378146 580580 604143
rect 580630 580816 580686 580825
rect 580630 580751 580686 580760
rect 580540 378140 580592 378146
rect 580540 378082 580592 378088
rect 580644 367062 580672 580751
rect 580722 557288 580778 557297
rect 580722 557223 580778 557232
rect 580632 367056 580684 367062
rect 580632 366998 580684 367004
rect 580736 362914 580764 557223
rect 580814 533896 580870 533905
rect 580814 533831 580870 533840
rect 580724 362908 580776 362914
rect 580724 362850 580776 362856
rect 580828 351898 580856 533831
rect 580906 510368 580962 510377
rect 580906 510303 580962 510312
rect 580816 351892 580868 351898
rect 580816 351834 580868 351840
rect 580920 346390 580948 510303
rect 580908 346384 580960 346390
rect 580908 346326 580960 346332
rect 580354 346080 580410 346089
rect 580354 346015 580410 346024
rect 580264 304972 580316 304978
rect 580264 304914 580316 304920
rect 580262 299160 580318 299169
rect 580262 299095 580318 299104
rect 392858 277672 392914 277681
rect 392858 277607 392914 277616
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 580184 274718 580212 275703
rect 392584 274712 392636 274718
rect 392584 274654 392636 274660
rect 580172 274712 580224 274718
rect 580172 274654 580224 274660
rect 152462 273592 152518 273601
rect 152462 273527 152518 273536
rect 3516 267776 3568 267782
rect 3516 267718 3568 267724
rect 3422 265704 3478 265713
rect 3422 265639 3478 265648
rect 3424 262268 3476 262274
rect 3424 262210 3476 262216
rect 3436 251297 3464 262210
rect 3422 251288 3478 251297
rect 3422 251223 3478 251232
rect 3424 249824 3476 249830
rect 3424 249766 3476 249772
rect 3148 208344 3200 208350
rect 3148 208286 3200 208292
rect 3160 208185 3188 208286
rect 3146 208176 3202 208185
rect 3146 208111 3202 208120
rect 3436 193905 3464 249766
rect 3528 237017 3556 267718
rect 3514 237008 3570 237017
rect 3514 236943 3570 236952
rect 3700 233300 3752 233306
rect 3700 233242 3752 233248
rect 3516 223576 3568 223582
rect 3516 223518 3568 223524
rect 3528 222601 3556 223518
rect 3514 222592 3570 222601
rect 3514 222527 3570 222536
rect 3608 216708 3660 216714
rect 3608 216650 3660 216656
rect 3516 200184 3568 200190
rect 3516 200126 3568 200132
rect 3422 193896 3478 193905
rect 3422 193831 3478 193840
rect 3424 182232 3476 182238
rect 3424 182174 3476 182180
rect 3056 180804 3108 180810
rect 3056 180746 3108 180752
rect 3068 179489 3096 180746
rect 3054 179480 3110 179489
rect 3054 179415 3110 179424
rect 3240 165572 3292 165578
rect 3240 165514 3292 165520
rect 3252 165073 3280 165514
rect 3238 165064 3294 165073
rect 3238 164999 3294 165008
rect 3332 136604 3384 136610
rect 3332 136546 3384 136552
rect 3344 136377 3372 136546
rect 3330 136368 3386 136377
rect 3330 136303 3386 136312
rect 3332 122800 3384 122806
rect 3332 122742 3384 122748
rect 3344 122097 3372 122742
rect 3330 122088 3386 122097
rect 3330 122023 3386 122032
rect 3056 80028 3108 80034
rect 3056 79970 3108 79976
rect 3068 78985 3096 79970
rect 3054 78976 3110 78985
rect 3054 78911 3110 78920
rect 3056 51060 3108 51066
rect 3056 51002 3108 51008
rect 3068 50153 3096 51002
rect 3054 50144 3110 50153
rect 3054 50079 3110 50088
rect 3436 21457 3464 182174
rect 3528 64569 3556 200126
rect 3620 107681 3648 216650
rect 3712 150793 3740 233242
rect 152476 223582 152504 273527
rect 391940 273216 391992 273222
rect 391940 273158 391992 273164
rect 391952 272377 391980 273158
rect 391938 272368 391994 272377
rect 391938 272303 391994 272312
rect 153106 268016 153162 268025
rect 153106 267951 153162 267960
rect 153120 267782 153148 267951
rect 153108 267776 153160 267782
rect 153108 267718 153160 267724
rect 392596 267073 392624 274654
rect 580276 273222 580304 299095
rect 580368 288386 580396 346015
rect 580356 288380 580408 288386
rect 580356 288322 580408 288328
rect 580264 273216 580316 273222
rect 580264 273158 580316 273164
rect 392582 267064 392638 267073
rect 392582 266999 392638 267008
rect 579802 263936 579858 263945
rect 579802 263871 579858 263880
rect 579816 263634 579844 263871
rect 391940 263628 391992 263634
rect 391940 263570 391992 263576
rect 579804 263628 579856 263634
rect 579804 263570 579856 263576
rect 153106 262304 153162 262313
rect 153106 262239 153108 262248
rect 153160 262239 153162 262248
rect 153108 262210 153160 262216
rect 391952 261905 391980 263570
rect 391938 261896 391994 261905
rect 391938 261831 391994 261840
rect 152646 256728 152702 256737
rect 152646 256663 152702 256672
rect 152554 245440 152610 245449
rect 152554 245375 152610 245384
rect 152464 223576 152516 223582
rect 152464 223518 152516 223524
rect 152568 208350 152596 245375
rect 152556 208344 152608 208350
rect 152556 208286 152608 208292
rect 152554 206000 152610 206009
rect 152554 205935 152610 205944
rect 152002 200288 152058 200297
rect 152002 200223 152058 200232
rect 152016 200190 152044 200223
rect 152004 200184 152056 200190
rect 152004 200126 152056 200132
rect 152278 189000 152334 189009
rect 152278 188935 152334 188944
rect 152292 180826 152320 188935
rect 152462 183424 152518 183433
rect 152462 183359 152518 183368
rect 152476 182238 152504 183359
rect 152464 182232 152516 182238
rect 152464 182174 152516 182180
rect 152292 180798 152504 180826
rect 122748 173732 122800 173738
rect 122748 173674 122800 173680
rect 118608 173664 118660 173670
rect 118608 173606 118660 173612
rect 111708 173596 111760 173602
rect 111708 173538 111760 173544
rect 35164 173528 35216 173534
rect 35164 173470 35216 173476
rect 29644 173460 29696 173466
rect 29644 173402 29696 173408
rect 19984 173392 20036 173398
rect 19984 173334 20036 173340
rect 18604 173256 18656 173262
rect 18604 173198 18656 173204
rect 10324 173188 10376 173194
rect 10324 173130 10376 173136
rect 3698 150784 3754 150793
rect 3698 150719 3754 150728
rect 3606 107672 3662 107681
rect 3606 107607 3662 107616
rect 3608 93832 3660 93838
rect 3608 93774 3660 93780
rect 3620 93265 3648 93774
rect 3606 93256 3662 93265
rect 3606 93191 3662 93200
rect 3514 64560 3570 64569
rect 3514 64495 3570 64504
rect 3516 35896 3568 35902
rect 3514 35864 3516 35873
rect 3568 35864 3570 35873
rect 3514 35799 3570 35808
rect 3422 21448 3478 21457
rect 3422 21383 3478 21392
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 7177 3464 8230
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 1676 4956 1728 4962
rect 1676 4898 1728 4904
rect 572 4820 624 4826
rect 572 4762 624 4768
rect 584 480 612 4762
rect 1688 480 1716 4898
rect 2872 4888 2924 4894
rect 2872 4830 2924 4836
rect 2884 480 2912 4830
rect 4080 480 4108 6122
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 5262 3360 5318 3369
rect 5262 3295 5318 3304
rect 5276 480 5304 3295
rect 6472 480 6500 3402
rect 7668 480 7696 4966
rect 8864 480 8892 6190
rect 10336 3466 10364 173130
rect 11704 158024 11756 158030
rect 11704 157966 11756 157972
rect 11242 3496 11298 3505
rect 10324 3460 10376 3466
rect 11242 3431 11298 3440
rect 10324 3402 10376 3408
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 10060 480 10088 2926
rect 11256 480 11284 3431
rect 11716 2990 11744 157966
rect 13636 10328 13688 10334
rect 13636 10270 13688 10276
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 12452 480 12480 5034
rect 13648 480 13676 10270
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 14844 480 14872 4082
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 16040 480 16068 3470
rect 17236 480 17264 5102
rect 18616 4146 18644 173198
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 19522 3632 19578 3641
rect 19522 3567 19578 3576
rect 18328 3324 18380 3330
rect 18328 3266 18380 3272
rect 18340 480 18368 3266
rect 19536 480 19564 3567
rect 19996 3534 20024 173334
rect 28264 173324 28316 173330
rect 28264 173266 28316 173272
rect 21364 162172 21416 162178
rect 21364 162114 21416 162120
rect 20718 3768 20774 3777
rect 20718 3703 20774 3712
rect 19984 3528 20036 3534
rect 19984 3470 20036 3476
rect 20732 480 20760 3703
rect 21376 3330 21404 162114
rect 23388 11756 23440 11762
rect 23388 11698 23440 11704
rect 21916 5228 21968 5234
rect 21916 5170 21968 5176
rect 21364 3324 21416 3330
rect 21364 3266 21416 3272
rect 21928 480 21956 5170
rect 23400 3482 23428 11698
rect 26700 5296 26752 5302
rect 26700 5238 26752 5244
rect 23124 3454 23428 3482
rect 25504 3528 25556 3534
rect 25504 3470 25556 3476
rect 23124 480 23152 3454
rect 24308 2984 24360 2990
rect 24308 2926 24360 2932
rect 24320 480 24348 2926
rect 25516 480 25544 3470
rect 26712 480 26740 5238
rect 27896 3256 27948 3262
rect 27896 3198 27948 3204
rect 27908 480 27936 3198
rect 28276 2990 28304 173266
rect 29656 3534 29684 173402
rect 32404 167680 32456 167686
rect 32404 167622 32456 167628
rect 31024 163532 31076 163538
rect 31024 163474 31076 163480
rect 30288 5364 30340 5370
rect 30288 5306 30340 5312
rect 29644 3528 29696 3534
rect 29644 3470 29696 3476
rect 29092 3460 29144 3466
rect 29092 3402 29144 3408
rect 28264 2984 28316 2990
rect 28264 2926 28316 2932
rect 29104 480 29132 3402
rect 30300 480 30328 5306
rect 31036 3262 31064 163474
rect 32416 3534 32444 167622
rect 33876 6316 33928 6322
rect 33876 6258 33928 6264
rect 31484 3528 31536 3534
rect 31484 3470 31536 3476
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 32680 3528 32732 3534
rect 32680 3470 32732 3476
rect 31024 3256 31076 3262
rect 31024 3198 31076 3204
rect 31496 480 31524 3470
rect 32692 480 32720 3470
rect 33888 480 33916 6258
rect 34980 3664 35032 3670
rect 34980 3606 35032 3612
rect 34992 480 35020 3606
rect 35176 3534 35204 173470
rect 36544 170400 36596 170406
rect 36544 170342 36596 170348
rect 36556 3670 36584 170342
rect 96528 169040 96580 169046
rect 96528 168982 96580 168988
rect 38568 166320 38620 166326
rect 38568 166262 38620 166268
rect 37372 6384 37424 6390
rect 37372 6326 37424 6332
rect 36544 3664 36596 3670
rect 36544 3606 36596 3612
rect 35164 3528 35216 3534
rect 35164 3470 35216 3476
rect 36176 3324 36228 3330
rect 36176 3266 36228 3272
rect 36188 480 36216 3266
rect 37384 480 37412 6326
rect 38580 480 38608 166262
rect 55128 160744 55180 160750
rect 55128 160686 55180 160692
rect 50988 156664 51040 156670
rect 50988 156606 51040 156612
rect 42708 155236 42760 155242
rect 42708 155178 42760 155184
rect 40960 6452 41012 6458
rect 40960 6394 41012 6400
rect 39764 3596 39816 3602
rect 39764 3538 39816 3544
rect 39776 480 39804 3538
rect 40972 480 41000 6394
rect 42720 3534 42748 155178
rect 46848 138712 46900 138718
rect 46848 138654 46900 138660
rect 44548 6520 44600 6526
rect 44548 6462 44600 6468
rect 43352 3664 43404 3670
rect 43352 3606 43404 3612
rect 42156 3528 42208 3534
rect 42156 3470 42208 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 42168 480 42196 3470
rect 43364 480 43392 3606
rect 44560 480 44588 6462
rect 46860 3398 46888 138654
rect 49332 7608 49384 7614
rect 49332 7550 49384 7556
rect 48136 5432 48188 5438
rect 48136 5374 48188 5380
rect 46940 3732 46992 3738
rect 46940 3674 46992 3680
rect 45744 3392 45796 3398
rect 45744 3334 45796 3340
rect 46848 3392 46900 3398
rect 46848 3334 46900 3340
rect 45756 480 45784 3334
rect 46952 480 46980 3674
rect 48148 480 48176 5374
rect 49344 480 49372 7550
rect 51000 3398 51028 156606
rect 52828 7676 52880 7682
rect 52828 7618 52880 7624
rect 51632 5500 51684 5506
rect 51632 5442 51684 5448
rect 50528 3392 50580 3398
rect 50528 3334 50580 3340
rect 50988 3392 51040 3398
rect 50988 3334 51040 3340
rect 50540 480 50568 3334
rect 51644 480 51672 5442
rect 52840 480 52868 7618
rect 55140 3398 55168 160686
rect 82728 153876 82780 153882
rect 82728 153818 82780 153824
rect 57888 137284 57940 137290
rect 57888 137226 57940 137232
rect 56416 7744 56468 7750
rect 56416 7686 56468 7692
rect 55220 4752 55272 4758
rect 55220 4694 55272 4700
rect 54024 3392 54076 3398
rect 54024 3334 54076 3340
rect 55128 3392 55180 3398
rect 55128 3334 55180 3340
rect 54036 480 54064 3334
rect 55232 480 55260 4694
rect 56428 480 56456 7686
rect 57900 626 57928 137226
rect 62028 134564 62080 134570
rect 62028 134506 62080 134512
rect 60004 7812 60056 7818
rect 60004 7754 60056 7760
rect 58808 4684 58860 4690
rect 58808 4626 58860 4632
rect 57624 598 57928 626
rect 57624 480 57652 598
rect 58820 480 58848 4626
rect 60016 480 60044 7754
rect 62040 3398 62068 134506
rect 77852 8152 77904 8158
rect 77852 8094 77904 8100
rect 74264 8084 74316 8090
rect 74264 8026 74316 8032
rect 70676 8016 70728 8022
rect 70676 7958 70728 7964
rect 67180 7948 67232 7954
rect 67180 7890 67232 7896
rect 63592 7880 63644 7886
rect 63592 7822 63644 7828
rect 62396 4616 62448 4622
rect 62396 4558 62448 4564
rect 61200 3392 61252 3398
rect 61200 3334 61252 3340
rect 62028 3392 62080 3398
rect 62028 3334 62080 3340
rect 61212 480 61240 3334
rect 62408 480 62436 4558
rect 63604 480 63632 7822
rect 65984 4548 66036 4554
rect 65984 4490 66036 4496
rect 64788 3800 64840 3806
rect 64788 3742 64840 3748
rect 64800 480 64828 3742
rect 65996 480 66024 4490
rect 67192 480 67220 7890
rect 69480 4480 69532 4486
rect 69480 4422 69532 4428
rect 68284 3868 68336 3874
rect 68284 3810 68336 3816
rect 68296 480 68324 3810
rect 69492 480 69520 4422
rect 70688 480 70716 7958
rect 73068 4412 73120 4418
rect 73068 4354 73120 4360
rect 71872 3936 71924 3942
rect 71872 3878 71924 3884
rect 71884 480 71912 3878
rect 73080 480 73108 4354
rect 74276 480 74304 8026
rect 76656 4344 76708 4350
rect 76656 4286 76708 4292
rect 75460 4004 75512 4010
rect 75460 3946 75512 3952
rect 75472 480 75500 3946
rect 76668 480 76696 4286
rect 77864 480 77892 8094
rect 80244 4276 80296 4282
rect 80244 4218 80296 4224
rect 79048 3256 79100 3262
rect 79048 3198 79100 3204
rect 79060 480 79088 3198
rect 80256 480 80284 4218
rect 82636 4072 82688 4078
rect 82636 4014 82688 4020
rect 81440 3392 81492 3398
rect 81440 3334 81492 3340
rect 81452 480 81480 3334
rect 82648 480 82676 4014
rect 82740 3398 82768 153818
rect 85488 152516 85540 152522
rect 85488 152458 85540 152464
rect 83832 6588 83884 6594
rect 83832 6530 83884 6536
rect 82728 3392 82780 3398
rect 82728 3334 82780 3340
rect 83844 480 83872 6530
rect 85500 3398 85528 152458
rect 89628 151088 89680 151094
rect 89628 151030 89680 151036
rect 87328 6656 87380 6662
rect 87328 6598 87380 6604
rect 84936 3392 84988 3398
rect 84936 3334 84988 3340
rect 85488 3392 85540 3398
rect 85488 3334 85540 3340
rect 84948 480 84976 3334
rect 86132 3256 86184 3262
rect 86132 3198 86184 3204
rect 86144 480 86172 3198
rect 87340 480 87368 6598
rect 89640 3398 89668 151030
rect 92388 149728 92440 149734
rect 92388 149670 92440 149676
rect 90916 6724 90968 6730
rect 90916 6666 90968 6672
rect 88524 3392 88576 3398
rect 88524 3334 88576 3340
rect 89628 3392 89680 3398
rect 89628 3334 89680 3340
rect 88536 480 88564 3334
rect 89904 3324 89956 3330
rect 89904 3266 89956 3272
rect 89916 1714 89944 3266
rect 89732 1686 89944 1714
rect 89732 480 89760 1686
rect 90928 480 90956 6666
rect 92400 3482 92428 149670
rect 94504 8220 94556 8226
rect 94504 8162 94556 8168
rect 92124 3454 92428 3482
rect 92124 480 92152 3454
rect 93308 3256 93360 3262
rect 93308 3198 93360 3204
rect 93320 480 93348 3198
rect 94516 480 94544 8162
rect 96540 3194 96568 168982
rect 99288 148368 99340 148374
rect 99288 148310 99340 148316
rect 98092 7540 98144 7546
rect 98092 7482 98144 7488
rect 95700 3188 95752 3194
rect 95700 3130 95752 3136
rect 96528 3188 96580 3194
rect 96528 3130 96580 3136
rect 95712 480 95740 3130
rect 96896 3052 96948 3058
rect 96896 2994 96948 3000
rect 96908 480 96936 2994
rect 98104 480 98132 7482
rect 99300 480 99328 148310
rect 103428 146940 103480 146946
rect 103428 146882 103480 146888
rect 101588 7472 101640 7478
rect 101588 7414 101640 7420
rect 100484 3120 100536 3126
rect 100484 3062 100536 3068
rect 100496 480 100524 3062
rect 101600 480 101628 7414
rect 103440 3194 103468 146882
rect 107568 145580 107620 145586
rect 107568 145522 107620 145528
rect 105176 7404 105228 7410
rect 105176 7346 105228 7352
rect 102784 3188 102836 3194
rect 102784 3130 102836 3136
rect 103428 3188 103480 3194
rect 103428 3130 103480 3136
rect 102796 480 102824 3130
rect 103980 2848 104032 2854
rect 103980 2790 104032 2796
rect 103992 480 104020 2790
rect 105188 480 105216 7346
rect 107580 3194 107608 145522
rect 110328 144220 110380 144226
rect 110328 144162 110380 144168
rect 108764 7336 108816 7342
rect 108764 7278 108816 7284
rect 106372 3188 106424 3194
rect 106372 3130 106424 3136
rect 107568 3188 107620 3194
rect 107568 3130 107620 3136
rect 106384 480 106412 3130
rect 107568 2848 107620 2854
rect 107568 2790 107620 2796
rect 107580 480 107608 2790
rect 108776 480 108804 7278
rect 110340 3482 110368 144162
rect 109972 3454 110368 3482
rect 109972 480 110000 3454
rect 111720 3194 111748 173538
rect 114468 171828 114520 171834
rect 114468 171770 114520 171776
rect 112352 7268 112404 7274
rect 112352 7210 112404 7216
rect 111156 3188 111208 3194
rect 111156 3130 111208 3136
rect 111708 3188 111760 3194
rect 111708 3130 111760 3136
rect 111168 480 111196 3130
rect 112364 480 112392 7210
rect 114480 2990 114508 171770
rect 117228 142860 117280 142866
rect 117228 142802 117280 142808
rect 115940 7200 115992 7206
rect 115940 7142 115992 7148
rect 113548 2984 113600 2990
rect 113548 2926 113600 2932
rect 114468 2984 114520 2990
rect 114468 2926 114520 2932
rect 113560 480 113588 2926
rect 114744 2916 114796 2922
rect 114744 2858 114796 2864
rect 114756 480 114784 2858
rect 115952 480 115980 7142
rect 117240 3482 117268 142802
rect 118620 3482 118648 173606
rect 121368 141432 121420 141438
rect 121368 141374 121420 141380
rect 119436 7132 119488 7138
rect 119436 7074 119488 7080
rect 117148 3454 117268 3482
rect 118252 3454 118648 3482
rect 117148 480 117176 3454
rect 118252 480 118280 3454
rect 119448 480 119476 7074
rect 121380 2990 121408 141374
rect 120632 2984 120684 2990
rect 120632 2926 120684 2932
rect 121368 2984 121420 2990
rect 121368 2926 121420 2932
rect 120644 480 120672 2926
rect 122760 2854 122788 173674
rect 126888 171896 126940 171902
rect 126888 171838 126940 171844
rect 125508 140072 125560 140078
rect 125508 140014 125560 140020
rect 123024 7064 123076 7070
rect 123024 7006 123076 7012
rect 121828 2848 121880 2854
rect 121828 2790 121880 2796
rect 122748 2848 122800 2854
rect 122748 2790 122800 2796
rect 121840 480 121868 2790
rect 123036 480 123064 7006
rect 125520 2854 125548 140014
rect 126900 3346 126928 171838
rect 131028 170468 131080 170474
rect 131028 170410 131080 170416
rect 128268 159384 128320 159390
rect 128268 159326 128320 159332
rect 126624 3318 126928 3346
rect 124220 2848 124272 2854
rect 124220 2790 124272 2796
rect 125508 2848 125560 2854
rect 125508 2790 125560 2796
rect 124232 480 124260 2790
rect 125416 2780 125468 2786
rect 125416 2722 125468 2728
rect 125428 480 125456 2722
rect 126624 480 126652 3318
rect 128280 2854 128308 159326
rect 129004 6792 129056 6798
rect 129004 6734 129056 6740
rect 127808 2848 127860 2854
rect 127808 2790 127860 2796
rect 128268 2848 128320 2854
rect 128268 2790 128320 2796
rect 127820 480 127848 2790
rect 129016 480 129044 6734
rect 131040 2854 131068 170410
rect 137928 169108 137980 169114
rect 137928 169050 137980 169056
rect 133788 166388 133840 166394
rect 133788 166330 133840 166336
rect 132408 160812 132460 160818
rect 132408 160754 132460 160760
rect 130200 2848 130252 2854
rect 130200 2790 130252 2796
rect 131028 2848 131080 2854
rect 131028 2790 131080 2796
rect 131396 2848 131448 2854
rect 131396 2790 131448 2796
rect 132316 2848 132368 2854
rect 132420 2836 132448 160754
rect 132592 6860 132644 6866
rect 132592 6802 132644 6808
rect 132368 2808 132448 2836
rect 132316 2790 132368 2796
rect 130212 480 130240 2790
rect 131408 480 131436 2790
rect 132604 480 132632 6802
rect 133800 480 133828 166330
rect 135168 17264 135220 17270
rect 135168 17206 135220 17212
rect 135180 626 135208 17206
rect 136088 6112 136140 6118
rect 136088 6054 136140 6060
rect 134904 598 135208 626
rect 134904 480 134932 598
rect 136100 480 136128 6054
rect 137940 610 137968 169050
rect 142068 167748 142120 167754
rect 142068 167690 142120 167696
rect 139308 156732 139360 156738
rect 139308 156674 139360 156680
rect 139320 610 139348 156674
rect 141976 22772 142028 22778
rect 141976 22714 142028 22720
rect 139676 6044 139728 6050
rect 139676 5986 139728 5992
rect 137284 604 137336 610
rect 137284 546 137336 552
rect 137928 604 137980 610
rect 137928 546 137980 552
rect 138480 604 138532 610
rect 138480 546 138532 552
rect 139308 604 139360 610
rect 139308 546 139360 552
rect 137296 480 137324 546
rect 138492 480 138520 546
rect 139688 480 139716 5986
rect 140872 4208 140924 4214
rect 140872 4150 140924 4156
rect 140884 480 140912 4150
rect 141988 3482 142016 22714
rect 142080 4214 142108 167690
rect 144828 164892 144880 164898
rect 144828 164834 144880 164840
rect 143264 5976 143316 5982
rect 143264 5918 143316 5924
rect 142068 4208 142120 4214
rect 142068 4150 142120 4156
rect 141988 3454 142108 3482
rect 142080 480 142108 3454
rect 143276 480 143304 5918
rect 144840 626 144868 164834
rect 148968 163600 149020 163606
rect 148968 163542 149020 163548
rect 146208 158092 146260 158098
rect 146208 158034 146260 158040
rect 144472 598 144868 626
rect 146220 610 146248 158034
rect 146852 5908 146904 5914
rect 146852 5850 146904 5856
rect 145656 604 145708 610
rect 144472 480 144500 598
rect 145656 546 145708 552
rect 146208 604 146260 610
rect 146208 546 146260 552
rect 145668 480 145696 546
rect 146864 480 146892 5850
rect 148980 610 149008 163542
rect 151728 162240 151780 162246
rect 151728 162182 151780 162188
rect 150348 155304 150400 155310
rect 150348 155246 150400 155252
rect 150360 610 150388 155246
rect 150440 5840 150492 5846
rect 150440 5782 150492 5788
rect 148048 604 148100 610
rect 148048 546 148100 552
rect 148968 604 149020 610
rect 148968 546 149020 552
rect 149244 604 149296 610
rect 149244 546 149296 552
rect 150348 604 150400 610
rect 150348 546 150400 552
rect 148060 480 148088 546
rect 149256 480 149284 546
rect 150452 480 150480 5782
rect 151740 610 151768 162182
rect 152476 8294 152504 180798
rect 152568 51066 152596 205935
rect 152660 180810 152688 256663
rect 391938 256592 391994 256601
rect 391938 256527 391994 256536
rect 391952 252550 391980 256527
rect 391940 252544 391992 252550
rect 391940 252486 391992 252492
rect 579804 252544 579856 252550
rect 579804 252486 579856 252492
rect 579816 252249 579844 252486
rect 579802 252240 579858 252249
rect 579802 252175 579858 252184
rect 392766 251288 392822 251297
rect 392766 251223 392822 251232
rect 153106 251016 153162 251025
rect 153106 250951 153162 250960
rect 153120 249830 153148 250951
rect 153108 249824 153160 249830
rect 153108 249766 153160 249772
rect 392674 245984 392730 245993
rect 392674 245919 392730 245928
rect 392582 240816 392638 240825
rect 392582 240751 392638 240760
rect 152922 239728 152978 239737
rect 152922 239663 152978 239672
rect 152738 222864 152794 222873
rect 152738 222799 152794 222808
rect 152648 180804 152700 180810
rect 152648 180746 152700 180752
rect 152646 177848 152702 177857
rect 152646 177783 152702 177792
rect 152556 51060 152608 51066
rect 152556 51002 152608 51008
rect 152660 35902 152688 177783
rect 152752 93838 152780 222799
rect 152830 194712 152886 194721
rect 152830 194647 152886 194656
rect 152740 93832 152792 93838
rect 152740 93774 152792 93780
rect 152844 80034 152872 194647
rect 152936 136610 152964 239663
rect 392490 235512 392546 235521
rect 392490 235447 392546 235456
rect 153106 234152 153162 234161
rect 153106 234087 153162 234096
rect 153120 233306 153148 234087
rect 153108 233300 153160 233306
rect 153108 233242 153160 233248
rect 153106 228576 153162 228585
rect 153106 228511 153162 228520
rect 153014 217288 153070 217297
rect 153014 217223 153070 217232
rect 153028 216714 153056 217223
rect 153016 216708 153068 216714
rect 153016 216650 153068 216656
rect 153014 211576 153070 211585
rect 153014 211511 153070 211520
rect 152924 136604 152976 136610
rect 152924 136546 152976 136552
rect 153028 122806 153056 211511
rect 153120 165578 153148 228511
rect 391938 209264 391994 209273
rect 391938 209199 391994 209208
rect 391952 208418 391980 209199
rect 391940 208412 391992 208418
rect 391940 208354 391992 208360
rect 392504 182170 392532 235447
rect 392596 205630 392624 240751
rect 392688 218006 392716 245919
rect 392780 229090 392808 251223
rect 393226 230208 393282 230217
rect 393226 230143 393282 230152
rect 392768 229084 392820 229090
rect 392768 229026 392820 229032
rect 393134 225040 393190 225049
rect 393134 224975 393190 224984
rect 393042 219736 393098 219745
rect 393042 219671 393098 219680
rect 392676 218000 392728 218006
rect 392676 217942 392728 217948
rect 392950 214432 393006 214441
rect 392950 214367 393006 214376
rect 392584 205624 392636 205630
rect 392584 205566 392636 205572
rect 392858 203960 392914 203969
rect 392858 203895 392914 203904
rect 392766 198656 392822 198665
rect 392766 198591 392822 198600
rect 392674 188184 392730 188193
rect 392674 188119 392730 188128
rect 392582 182880 392638 182889
rect 392582 182815 392638 182824
rect 392492 182164 392544 182170
rect 392492 182106 392544 182112
rect 391938 177712 391994 177721
rect 391938 177647 391994 177656
rect 391952 176730 391980 177647
rect 391940 176724 391992 176730
rect 391940 176666 391992 176672
rect 159100 175222 159482 175250
rect 166276 175222 166658 175250
rect 184492 175222 184874 175250
rect 185412 175222 185886 175250
rect 196452 175222 196834 175250
rect 197924 175222 198306 175250
rect 206572 175222 206954 175250
rect 217060 175222 217442 175250
rect 219912 175222 220386 175250
rect 224236 175222 224618 175250
rect 227088 175222 227562 175250
rect 229480 175222 229954 175250
rect 242452 175222 242834 175250
rect 256896 175222 257186 175250
rect 274022 175222 274404 175250
rect 282118 175222 282500 175250
rect 304198 175222 304580 175250
rect 309902 175222 310284 175250
rect 319470 175222 319852 175250
rect 320942 175222 321324 175250
rect 341550 175222 341932 175250
rect 342930 175222 343404 175250
rect 154684 175086 155250 175114
rect 155328 175086 155710 175114
rect 156064 175086 156170 175114
rect 156248 175086 156630 175114
rect 156892 175086 157090 175114
rect 154580 171080 154632 171086
rect 154580 171022 154632 171028
rect 153108 165572 153160 165578
rect 153108 165514 153160 165520
rect 153016 122800 153068 122806
rect 153016 122742 153068 122748
rect 152832 80028 152884 80034
rect 152832 79970 152884 79976
rect 152648 35896 152700 35902
rect 152648 35838 152700 35844
rect 153108 24132 153160 24138
rect 153108 24074 153160 24080
rect 152464 8288 152516 8294
rect 152464 8230 152516 8236
rect 153120 626 153148 24074
rect 153936 5772 153988 5778
rect 153936 5714 153988 5720
rect 151544 604 151596 610
rect 151544 546 151596 552
rect 151728 604 151780 610
rect 151728 546 151780 552
rect 152752 598 153148 626
rect 151556 480 151584 546
rect 152752 480 152780 598
rect 153948 480 153976 5714
rect 154592 4962 154620 171022
rect 154580 4956 154632 4962
rect 154580 4898 154632 4904
rect 154684 4826 154712 175086
rect 155328 171086 155356 175086
rect 155316 171080 155368 171086
rect 155316 171022 155368 171028
rect 156064 4894 156092 175086
rect 156248 171034 156276 175086
rect 156156 171006 156276 171034
rect 156156 6186 156184 171006
rect 156892 167074 156920 175086
rect 157628 173194 157656 175100
rect 157812 175086 158102 175114
rect 158272 175086 158562 175114
rect 158916 175086 159022 175114
rect 157616 173188 157668 173194
rect 157616 173130 157668 173136
rect 157432 168360 157484 168366
rect 157432 168302 157484 168308
rect 156236 167068 156288 167074
rect 156236 167010 156288 167016
rect 156880 167068 156932 167074
rect 156880 167010 156932 167016
rect 156248 157298 156276 167010
rect 156248 157270 156460 157298
rect 156432 147694 156460 157270
rect 156236 147688 156288 147694
rect 156236 147630 156288 147636
rect 156420 147688 156472 147694
rect 156420 147630 156472 147636
rect 156248 137986 156276 147630
rect 156248 137958 156460 137986
rect 156432 128382 156460 137958
rect 156236 128376 156288 128382
rect 156236 128318 156288 128324
rect 156420 128376 156472 128382
rect 156420 128318 156472 128324
rect 156248 118674 156276 128318
rect 156248 118646 156460 118674
rect 156432 109070 156460 118646
rect 156236 109064 156288 109070
rect 156236 109006 156288 109012
rect 156420 109064 156472 109070
rect 156420 109006 156472 109012
rect 156248 99362 156276 109006
rect 156248 99334 156460 99362
rect 156432 89758 156460 99334
rect 156236 89752 156288 89758
rect 156236 89694 156288 89700
rect 156420 89752 156472 89758
rect 156420 89694 156472 89700
rect 156248 80050 156276 89694
rect 156248 80022 156460 80050
rect 156432 50946 156460 80022
rect 156340 50918 156460 50946
rect 156340 41426 156368 50918
rect 156340 41398 156460 41426
rect 156432 31770 156460 41398
rect 156248 31742 156460 31770
rect 156248 22098 156276 31742
rect 157248 25560 157300 25566
rect 157248 25502 157300 25508
rect 156236 22092 156288 22098
rect 156236 22034 156288 22040
rect 156420 22092 156472 22098
rect 156420 22034 156472 22040
rect 156432 19310 156460 22034
rect 156420 19304 156472 19310
rect 156420 19246 156472 19252
rect 156420 12436 156472 12442
rect 156420 12378 156472 12384
rect 156144 6180 156196 6186
rect 156144 6122 156196 6128
rect 156052 4888 156104 4894
rect 156052 4830 156104 4836
rect 154672 4820 154724 4826
rect 154672 4762 154724 4768
rect 155132 4820 155184 4826
rect 155132 4762 155184 4768
rect 155144 480 155172 4762
rect 156432 3369 156460 12378
rect 156418 3360 156474 3369
rect 156418 3295 156474 3304
rect 157260 610 157288 25502
rect 157444 6254 157472 168302
rect 157812 154601 157840 175086
rect 158272 168366 158300 175086
rect 158260 168360 158312 168366
rect 158260 168302 158312 168308
rect 158812 168360 158864 168366
rect 158812 168302 158864 168308
rect 157614 154592 157670 154601
rect 157614 154527 157670 154536
rect 157798 154592 157854 154601
rect 157798 154527 157854 154536
rect 157628 145081 157656 154527
rect 157614 145072 157670 145081
rect 157614 145007 157670 145016
rect 157614 144936 157670 144945
rect 157614 144871 157670 144880
rect 157628 138106 157656 144871
rect 157616 138100 157668 138106
rect 157616 138042 157668 138048
rect 157616 137964 157668 137970
rect 157616 137906 157668 137912
rect 157628 133906 157656 137906
rect 157628 133890 157840 133906
rect 157628 133884 157852 133890
rect 157628 133878 157800 133884
rect 157800 133826 157852 133832
rect 157812 133795 157840 133826
rect 157616 124228 157668 124234
rect 157616 124170 157668 124176
rect 157628 109070 157656 124170
rect 157616 109064 157668 109070
rect 157616 109006 157668 109012
rect 157708 108996 157760 109002
rect 157708 108938 157760 108944
rect 157536 99414 157564 99445
rect 157720 99414 157748 108938
rect 157524 99408 157576 99414
rect 157708 99408 157760 99414
rect 157576 99356 157656 99362
rect 157524 99350 157656 99356
rect 157708 99350 157760 99356
rect 157536 99334 157656 99350
rect 157628 89758 157656 99334
rect 157616 89752 157668 89758
rect 157616 89694 157668 89700
rect 157708 89616 157760 89622
rect 157708 89558 157760 89564
rect 157536 80102 157564 80133
rect 157720 80102 157748 89558
rect 157524 80096 157576 80102
rect 157708 80096 157760 80102
rect 157576 80044 157656 80050
rect 157524 80038 157656 80044
rect 157708 80038 157760 80044
rect 157536 80022 157656 80038
rect 157628 70446 157656 80022
rect 158720 75948 158772 75954
rect 158720 75890 158772 75896
rect 157616 70440 157668 70446
rect 157616 70382 157668 70388
rect 157708 70304 157760 70310
rect 157708 70246 157760 70252
rect 157720 60738 157748 70246
rect 158732 67697 158760 75890
rect 158718 67688 158774 67697
rect 158718 67623 158774 67632
rect 157536 60710 157748 60738
rect 157536 60602 157564 60710
rect 157536 60574 157656 60602
rect 157628 53122 157656 60574
rect 157536 53094 157656 53122
rect 157536 50946 157564 53094
rect 157536 50918 157748 50946
rect 157720 41426 157748 50918
rect 157536 41398 157748 41426
rect 157536 41290 157564 41398
rect 157536 41262 157656 41290
rect 157628 21978 157656 41262
rect 157628 21950 157748 21978
rect 157432 6248 157484 6254
rect 157432 6190 157484 6196
rect 157524 6180 157576 6186
rect 157524 6122 157576 6128
rect 156328 604 156380 610
rect 156328 546 156380 552
rect 157248 604 157300 610
rect 157248 546 157300 552
rect 156340 480 156368 546
rect 157536 480 157564 6122
rect 157720 5030 157748 21950
rect 158824 5098 158852 168302
rect 158916 158030 158944 175086
rect 159100 169182 159128 175222
rect 159744 175086 160034 175114
rect 160204 175086 160494 175114
rect 159088 169176 159140 169182
rect 159088 169118 159140 169124
rect 159272 169176 159324 169182
rect 159272 169118 159324 169124
rect 159284 164257 159312 169118
rect 159744 168366 159772 175086
rect 159732 168360 159784 168366
rect 159732 168302 159784 168308
rect 159086 164248 159142 164257
rect 159086 164183 159142 164192
rect 159270 164248 159326 164257
rect 159270 164183 159326 164192
rect 159100 159338 159128 164183
rect 159008 159310 159128 159338
rect 158904 158024 158956 158030
rect 158904 157966 158956 157972
rect 159008 145081 159036 159310
rect 158994 145072 159050 145081
rect 158994 145007 159050 145016
rect 158994 144936 159050 144945
rect 158994 144871 159050 144880
rect 159008 143546 159036 144871
rect 158996 143540 159048 143546
rect 158996 143482 159048 143488
rect 159088 131028 159140 131034
rect 159088 130970 159140 130976
rect 159100 122806 159128 130970
rect 159088 122800 159140 122806
rect 159088 122742 159140 122748
rect 158904 113212 158956 113218
rect 158904 113154 158956 113160
rect 158916 113082 158944 113154
rect 158904 113076 158956 113082
rect 158904 113018 158956 113024
rect 159088 103556 159140 103562
rect 159088 103498 159140 103504
rect 159100 95266 159128 103498
rect 158904 95260 158956 95266
rect 158904 95202 158956 95208
rect 159088 95260 159140 95266
rect 159088 95202 159140 95208
rect 158916 95130 158944 95202
rect 158904 95124 158956 95130
rect 158904 95066 158956 95072
rect 158996 85604 159048 85610
rect 158996 85546 159048 85552
rect 159008 85490 159036 85546
rect 158916 85462 159036 85490
rect 158916 75954 158944 85462
rect 158904 75948 158956 75954
rect 158904 75890 158956 75896
rect 158994 67688 159050 67697
rect 158994 67623 159050 67632
rect 159008 66230 159036 67623
rect 158996 66224 159048 66230
rect 158996 66166 159048 66172
rect 158996 56636 159048 56642
rect 158996 56578 159048 56584
rect 159008 48346 159036 56578
rect 158996 48340 159048 48346
rect 158996 48282 159048 48288
rect 158904 48272 158956 48278
rect 158904 48214 158956 48220
rect 158916 46918 158944 48214
rect 158904 46912 158956 46918
rect 158904 46854 158956 46860
rect 159916 29640 159968 29646
rect 159916 29582 159968 29588
rect 158904 29096 158956 29102
rect 158904 29038 158956 29044
rect 158916 27606 158944 29038
rect 158904 27600 158956 27606
rect 158904 27542 158956 27548
rect 158904 19236 158956 19242
rect 158904 19178 158956 19184
rect 158916 9722 158944 19178
rect 158904 9716 158956 9722
rect 158904 9658 158956 9664
rect 158996 9716 159048 9722
rect 158996 9658 159048 9664
rect 158812 5092 158864 5098
rect 158812 5034 158864 5040
rect 157708 5024 157760 5030
rect 157708 4966 157760 4972
rect 158720 4888 158772 4894
rect 158720 4830 158772 4836
rect 158732 480 158760 4830
rect 159008 3505 159036 9658
rect 158994 3496 159050 3505
rect 158994 3431 159050 3440
rect 159928 480 159956 29582
rect 160204 10334 160232 175086
rect 160940 173262 160968 175100
rect 161400 173398 161428 175100
rect 161492 175086 161874 175114
rect 162044 175086 162426 175114
rect 161388 173392 161440 173398
rect 161388 173334 161440 173340
rect 160928 173256 160980 173262
rect 160928 173198 160980 173204
rect 160192 10328 160244 10334
rect 160192 10270 160244 10276
rect 161112 6248 161164 6254
rect 161112 6190 161164 6196
rect 161124 480 161152 6190
rect 161492 5166 161520 175086
rect 162044 167056 162072 175086
rect 161584 167028 162072 167056
rect 161584 162178 161612 167028
rect 161572 162172 161624 162178
rect 161572 162114 161624 162120
rect 162308 8968 162360 8974
rect 162308 8910 162360 8916
rect 161480 5160 161532 5166
rect 161480 5102 161532 5108
rect 162320 480 162348 8910
rect 162872 3641 162900 175100
rect 162964 175086 163346 175114
rect 163516 175086 163806 175114
rect 164266 175086 164372 175114
rect 162964 3777 162992 175086
rect 163516 172514 163544 175086
rect 163504 172508 163556 172514
rect 163504 172450 163556 172456
rect 163044 162920 163096 162926
rect 163096 162868 163176 162874
rect 163044 162862 163176 162868
rect 163056 162858 163176 162862
rect 163056 162852 163188 162858
rect 163056 162846 163136 162852
rect 163136 162794 163188 162800
rect 163320 162852 163372 162858
rect 163320 162794 163372 162800
rect 163332 161430 163360 162794
rect 163320 161424 163372 161430
rect 163320 161366 163372 161372
rect 163044 151836 163096 151842
rect 163044 151778 163096 151784
rect 163056 143585 163084 151778
rect 163042 143576 163098 143585
rect 163042 143511 163098 143520
rect 163226 143576 163282 143585
rect 163226 143511 163228 143520
rect 163280 143511 163282 143520
rect 163228 143482 163280 143488
rect 163136 128308 163188 128314
rect 163136 128250 163188 128256
rect 163148 125610 163176 128250
rect 163148 125582 163268 125610
rect 163056 118726 163084 118757
rect 163240 118726 163268 125582
rect 163044 118720 163096 118726
rect 163228 118720 163280 118726
rect 163096 118668 163176 118674
rect 163044 118662 163176 118668
rect 163228 118662 163280 118668
rect 163056 118646 163176 118662
rect 163148 115938 163176 118646
rect 163136 115932 163188 115938
rect 163136 115874 163188 115880
rect 163136 108996 163188 109002
rect 163136 108938 163188 108944
rect 163148 106298 163176 108938
rect 163148 106270 163268 106298
rect 163056 99414 163084 99445
rect 163240 99414 163268 106270
rect 163044 99408 163096 99414
rect 163228 99408 163280 99414
rect 163096 99356 163176 99362
rect 163044 99350 163176 99356
rect 163228 99350 163280 99356
rect 163056 99334 163176 99350
rect 163148 96626 163176 99334
rect 163136 96620 163188 96626
rect 163136 96562 163188 96568
rect 163136 89684 163188 89690
rect 163136 89626 163188 89632
rect 163148 86986 163176 89626
rect 163148 86958 163268 86986
rect 163056 80102 163084 80133
rect 163240 80102 163268 86958
rect 163044 80096 163096 80102
rect 163228 80096 163280 80102
rect 163096 80044 163176 80050
rect 163044 80038 163176 80044
rect 163228 80038 163280 80044
rect 163056 80022 163176 80038
rect 163148 70446 163176 80022
rect 163136 70440 163188 70446
rect 163136 70382 163188 70388
rect 163228 70304 163280 70310
rect 163228 70246 163280 70252
rect 163240 60738 163268 70246
rect 163056 60710 163268 60738
rect 163056 60602 163084 60710
rect 163056 60574 163176 60602
rect 163148 53122 163176 60574
rect 163056 53094 163176 53122
rect 163056 50946 163084 53094
rect 163056 50918 163268 50946
rect 163240 41426 163268 50918
rect 163056 41398 163268 41426
rect 163056 41290 163084 41398
rect 163056 41262 163176 41290
rect 163148 38622 163176 41262
rect 163136 38616 163188 38622
rect 163136 38558 163188 38564
rect 163228 29028 163280 29034
rect 163228 28970 163280 28976
rect 163240 22114 163268 28970
rect 163056 22086 163268 22114
rect 163056 21978 163084 22086
rect 163056 21950 163176 21978
rect 163148 5234 163176 21950
rect 164344 11762 164372 175086
rect 164804 173330 164832 175100
rect 165264 173466 165292 175100
rect 165252 173460 165304 173466
rect 165252 173402 165304 173408
rect 164792 173324 164844 173330
rect 164792 173266 164844 173272
rect 164332 11756 164384 11762
rect 164332 11698 164384 11704
rect 164700 5704 164752 5710
rect 164700 5646 164752 5652
rect 163136 5228 163188 5234
rect 163136 5170 163188 5176
rect 163504 4956 163556 4962
rect 163504 4898 163556 4904
rect 162950 3768 163006 3777
rect 162950 3703 163006 3712
rect 162858 3632 162914 3641
rect 162858 3567 162914 3576
rect 163516 480 163544 4898
rect 164712 480 164740 5646
rect 165724 5302 165752 175100
rect 165816 175086 166198 175114
rect 165816 163538 165844 175086
rect 166276 167056 166304 175222
rect 165908 167028 166304 167056
rect 165804 163532 165856 163538
rect 165804 163474 165856 163480
rect 165908 162194 165936 167028
rect 165816 162166 165936 162194
rect 165816 157298 165844 162166
rect 165816 157270 165936 157298
rect 165908 12458 165936 157270
rect 165816 12430 165936 12458
rect 165712 5296 165764 5302
rect 165712 5238 165764 5244
rect 165816 3670 165844 12430
rect 165896 10328 165948 10334
rect 165896 10270 165948 10276
rect 165804 3664 165856 3670
rect 165804 3606 165856 3612
rect 165908 480 165936 10270
rect 167196 5370 167224 175100
rect 167656 167686 167684 175100
rect 168116 173534 168144 175100
rect 168484 175086 168590 175114
rect 168104 173528 168156 173534
rect 168104 173470 168156 173476
rect 167644 167680 167696 167686
rect 167644 167622 167696 167628
rect 168380 164212 168432 164218
rect 168380 164154 168432 164160
rect 168392 154601 168420 164154
rect 168378 154592 168434 154601
rect 168378 154527 168434 154536
rect 168380 143540 168432 143546
rect 168380 143482 168432 143488
rect 168392 133929 168420 143482
rect 168378 133920 168434 133929
rect 168378 133855 168434 133864
rect 168484 6322 168512 175086
rect 169036 170406 169064 175100
rect 169220 175086 169602 175114
rect 169864 175086 170062 175114
rect 170324 175086 170522 175114
rect 170600 175086 170982 175114
rect 171244 175086 171534 175114
rect 171796 175086 171994 175114
rect 172072 175086 172454 175114
rect 172532 175086 172914 175114
rect 173084 175086 173374 175114
rect 169024 170400 169076 170406
rect 169024 170342 169076 170348
rect 169220 170218 169248 175086
rect 169760 171080 169812 171086
rect 169760 171022 169812 171028
rect 168668 170190 169248 170218
rect 168668 164218 168696 170190
rect 168656 164212 168708 164218
rect 168656 164154 168708 164160
rect 168562 154592 168618 154601
rect 168562 154527 168618 154536
rect 168576 147694 168604 154527
rect 168564 147688 168616 147694
rect 168564 147630 168616 147636
rect 168656 147620 168708 147626
rect 168656 147562 168708 147568
rect 168668 143546 168696 147562
rect 168656 143540 168708 143546
rect 168656 143482 168708 143488
rect 168562 133920 168618 133929
rect 168562 133855 168618 133864
rect 168576 124114 168604 133855
rect 168576 124086 168696 124114
rect 168668 114578 168696 124086
rect 168564 114572 168616 114578
rect 168564 114514 168616 114520
rect 168656 114572 168708 114578
rect 168656 114514 168708 114520
rect 168576 104802 168604 114514
rect 168576 104774 168696 104802
rect 168668 95266 168696 104774
rect 168564 95260 168616 95266
rect 168564 95202 168616 95208
rect 168656 95260 168708 95266
rect 168656 95202 168708 95208
rect 168576 77194 168604 95202
rect 168576 77166 168696 77194
rect 168668 67658 168696 77166
rect 168564 67652 168616 67658
rect 168564 67594 168616 67600
rect 168656 67652 168708 67658
rect 168656 67594 168708 67600
rect 168576 67538 168604 67594
rect 168576 67510 168696 67538
rect 168668 58002 168696 67510
rect 168564 57996 168616 58002
rect 168564 57938 168616 57944
rect 168656 57996 168708 58002
rect 168656 57938 168708 57944
rect 168576 48226 168604 57938
rect 168576 48198 168696 48226
rect 168668 38690 168696 48198
rect 168564 38684 168616 38690
rect 168564 38626 168616 38632
rect 168656 38684 168708 38690
rect 168656 38626 168708 38632
rect 168576 28914 168604 38626
rect 168576 28886 168788 28914
rect 168472 6316 168524 6322
rect 168472 6258 168524 6264
rect 168196 5636 168248 5642
rect 168196 5578 168248 5584
rect 167184 5364 167236 5370
rect 167184 5306 167236 5312
rect 167092 5024 167144 5030
rect 167092 4966 167144 4972
rect 167104 480 167132 4966
rect 168208 480 168236 5578
rect 168760 3534 168788 28886
rect 169392 11756 169444 11762
rect 169392 11698 169444 11704
rect 168748 3528 168800 3534
rect 168748 3470 168800 3476
rect 169404 480 169432 11698
rect 169772 3602 169800 171022
rect 169864 6390 169892 175086
rect 170324 171034 170352 175086
rect 170600 171086 170628 175086
rect 169956 171006 170352 171034
rect 170588 171080 170640 171086
rect 170588 171022 170640 171028
rect 171140 171080 171192 171086
rect 171140 171022 171192 171028
rect 169956 166326 169984 171006
rect 169944 166320 169996 166326
rect 169944 166262 169996 166268
rect 169852 6384 169904 6390
rect 169852 6326 169904 6332
rect 170588 5092 170640 5098
rect 170588 5034 170640 5040
rect 169760 3596 169812 3602
rect 169760 3538 169812 3544
rect 170600 480 170628 5034
rect 171152 3466 171180 171022
rect 171244 6458 171272 175086
rect 171796 171034 171824 175086
rect 172072 171086 172100 175086
rect 171428 171006 171824 171034
rect 172060 171080 172112 171086
rect 172060 171022 172112 171028
rect 171428 155242 171456 171006
rect 172428 164212 172480 164218
rect 172428 164154 172480 164160
rect 171416 155236 171468 155242
rect 171416 155178 171468 155184
rect 172440 154601 172468 164154
rect 172426 154592 172482 154601
rect 172426 154527 172482 154536
rect 172532 6526 172560 175086
rect 173084 171034 173112 175086
rect 172716 171006 173112 171034
rect 172716 164218 172744 171006
rect 172704 164212 172756 164218
rect 172704 164154 172756 164160
rect 172610 154592 172666 154601
rect 172610 154527 172666 154536
rect 172624 138718 172652 154527
rect 172612 138712 172664 138718
rect 172612 138654 172664 138660
rect 173808 18624 173860 18630
rect 173808 18566 173860 18572
rect 172520 6520 172572 6526
rect 172520 6462 172572 6468
rect 171232 6452 171284 6458
rect 171232 6394 171284 6400
rect 171784 6316 171836 6322
rect 171784 6258 171836 6264
rect 171140 3460 171192 3466
rect 171140 3402 171192 3408
rect 171796 480 171824 6258
rect 173820 3874 173848 18566
rect 172980 3868 173032 3874
rect 172980 3810 173032 3816
rect 173808 3868 173860 3874
rect 173808 3810 173860 3816
rect 172992 480 173020 3810
rect 173912 3738 173940 175100
rect 174004 175086 174386 175114
rect 174556 175086 174846 175114
rect 175306 175086 175504 175114
rect 174004 5438 174032 175086
rect 174556 165374 174584 175086
rect 175372 171080 175424 171086
rect 175372 171022 175424 171028
rect 175280 171012 175332 171018
rect 175280 170954 175332 170960
rect 174084 165368 174136 165374
rect 174084 165310 174136 165316
rect 174544 165368 174596 165374
rect 174544 165310 174596 165316
rect 174096 162858 174124 165310
rect 174084 162852 174136 162858
rect 174084 162794 174136 162800
rect 174268 162852 174320 162858
rect 174268 162794 174320 162800
rect 174280 128382 174308 162794
rect 174084 128376 174136 128382
rect 174268 128376 174320 128382
rect 174136 128324 174216 128330
rect 174084 128318 174216 128324
rect 174268 128318 174320 128324
rect 174096 128302 174216 128318
rect 174188 118726 174216 128302
rect 174176 118720 174228 118726
rect 174176 118662 174228 118668
rect 174268 118652 174320 118658
rect 174268 118594 174320 118600
rect 174280 109070 174308 118594
rect 174084 109064 174136 109070
rect 174268 109064 174320 109070
rect 174136 109012 174216 109018
rect 174084 109006 174216 109012
rect 174268 109006 174320 109012
rect 174096 108990 174216 109006
rect 174188 104854 174216 108990
rect 174176 104848 174228 104854
rect 174176 104790 174228 104796
rect 174268 95260 174320 95266
rect 174268 95202 174320 95208
rect 174280 89758 174308 95202
rect 174084 89752 174136 89758
rect 174268 89752 174320 89758
rect 174136 89700 174216 89706
rect 174084 89694 174216 89700
rect 174268 89694 174320 89700
rect 174096 89678 174216 89694
rect 174188 85542 174216 89678
rect 174176 85536 174228 85542
rect 174176 85478 174228 85484
rect 174268 75948 174320 75954
rect 174268 75890 174320 75896
rect 174280 66298 174308 75890
rect 174176 66292 174228 66298
rect 174176 66234 174228 66240
rect 174268 66292 174320 66298
rect 174268 66234 174320 66240
rect 174188 60738 174216 66234
rect 174188 60710 174308 60738
rect 174280 50946 174308 60710
rect 174188 50918 174308 50946
rect 174188 41426 174216 50918
rect 174188 41398 174308 41426
rect 174280 29102 174308 41398
rect 174268 29096 174320 29102
rect 174268 29038 174320 29044
rect 174176 29028 174228 29034
rect 174176 28970 174228 28976
rect 174188 22114 174216 28970
rect 174188 22086 174308 22114
rect 174280 12458 174308 22086
rect 174096 12430 174308 12458
rect 174096 7614 174124 12430
rect 174084 7608 174136 7614
rect 174084 7550 174136 7556
rect 175292 5506 175320 170954
rect 175384 7682 175412 171022
rect 175476 156670 175504 175086
rect 175568 175086 175766 175114
rect 175936 175086 176318 175114
rect 176778 175086 176884 175114
rect 175568 171018 175596 175086
rect 175936 171086 175964 175086
rect 175924 171080 175976 171086
rect 175924 171022 175976 171028
rect 176660 171080 176712 171086
rect 176660 171022 176712 171028
rect 175556 171012 175608 171018
rect 175556 170954 175608 170960
rect 175464 156664 175516 156670
rect 175464 156606 175516 156612
rect 176568 13116 176620 13122
rect 176568 13058 176620 13064
rect 175372 7676 175424 7682
rect 175372 7618 175424 7624
rect 175372 6384 175424 6390
rect 175372 6326 175424 6332
rect 175280 5500 175332 5506
rect 175280 5442 175332 5448
rect 173992 5432 174044 5438
rect 173992 5374 174044 5380
rect 174176 5160 174228 5166
rect 174176 5102 174228 5108
rect 173900 3732 173952 3738
rect 173900 3674 173952 3680
rect 174188 480 174216 5102
rect 175384 480 175412 6326
rect 176580 480 176608 13058
rect 176672 4758 176700 171022
rect 176752 171012 176804 171018
rect 176752 170954 176804 170960
rect 176764 7750 176792 170954
rect 176856 160750 176884 175086
rect 177132 175086 177238 175114
rect 177408 175086 177698 175114
rect 178158 175086 178264 175114
rect 177132 171086 177160 175086
rect 177120 171080 177172 171086
rect 177120 171022 177172 171028
rect 177408 171018 177436 175086
rect 178040 171080 178092 171086
rect 178040 171022 178092 171028
rect 177396 171012 177448 171018
rect 177396 170954 177448 170960
rect 176844 160744 176896 160750
rect 176844 160686 176896 160692
rect 176752 7744 176804 7750
rect 176752 7686 176804 7692
rect 177764 5228 177816 5234
rect 177764 5170 177816 5176
rect 176660 4752 176712 4758
rect 176660 4694 176712 4700
rect 177776 480 177804 5170
rect 178052 4690 178080 171022
rect 178132 167680 178184 167686
rect 178132 167622 178184 167628
rect 178144 7818 178172 167622
rect 178236 137290 178264 175086
rect 178328 175086 178710 175114
rect 178880 175086 179170 175114
rect 179524 175086 179630 175114
rect 179892 175086 180090 175114
rect 180168 175086 180550 175114
rect 180812 175086 181102 175114
rect 181180 175086 181562 175114
rect 181732 175086 182022 175114
rect 182192 175086 182482 175114
rect 182560 175086 182942 175114
rect 183204 175086 183494 175114
rect 183572 175086 183954 175114
rect 184032 175086 184414 175114
rect 178328 171086 178356 175086
rect 178316 171080 178368 171086
rect 178316 171022 178368 171028
rect 178880 167686 178908 175086
rect 179524 172553 179552 175086
rect 179510 172544 179566 172553
rect 179510 172479 179566 172488
rect 179694 172544 179750 172553
rect 179694 172479 179750 172488
rect 179420 171080 179472 171086
rect 179420 171022 179472 171028
rect 178868 167680 178920 167686
rect 178868 167622 178920 167628
rect 178224 137284 178276 137290
rect 178224 137226 178276 137232
rect 178132 7812 178184 7818
rect 178132 7754 178184 7760
rect 178960 6452 179012 6458
rect 178960 6394 179012 6400
rect 178040 4684 178092 4690
rect 178040 4626 178092 4632
rect 178972 480 179000 6394
rect 179432 4622 179460 171022
rect 179512 171012 179564 171018
rect 179512 170954 179564 170960
rect 179524 7886 179552 170954
rect 179708 167668 179736 172479
rect 179892 171086 179920 175086
rect 179880 171080 179932 171086
rect 179880 171022 179932 171028
rect 180168 171018 180196 175086
rect 180156 171012 180208 171018
rect 180156 170954 180208 170960
rect 179708 167640 179920 167668
rect 179892 153241 179920 167640
rect 179694 153232 179750 153241
rect 179616 153190 179694 153218
rect 179616 143546 179644 153190
rect 179694 153167 179750 153176
rect 179878 153232 179934 153241
rect 179878 153167 179934 153176
rect 179604 143540 179656 143546
rect 179604 143482 179656 143488
rect 180708 19984 180760 19990
rect 180708 19926 180760 19932
rect 179512 7880 179564 7886
rect 179512 7822 179564 7828
rect 179420 4616 179472 4622
rect 179420 4558 179472 4564
rect 180720 4010 180748 19926
rect 180156 4004 180208 4010
rect 180156 3946 180208 3952
rect 180708 4004 180760 4010
rect 180708 3946 180760 3952
rect 180168 480 180196 3946
rect 180812 3738 180840 175086
rect 181180 171068 181208 175086
rect 180904 171040 181208 171068
rect 180904 4554 180932 171040
rect 181732 164286 181760 175086
rect 181168 164280 181220 164286
rect 181168 164222 181220 164228
rect 181720 164280 181772 164286
rect 181720 164222 181772 164228
rect 181180 162858 181208 164222
rect 181168 162852 181220 162858
rect 181168 162794 181220 162800
rect 181168 145036 181220 145042
rect 181168 144978 181220 144984
rect 181180 143546 181208 144978
rect 181168 143540 181220 143546
rect 181168 143482 181220 143488
rect 181076 134020 181128 134026
rect 181076 133962 181128 133968
rect 181088 133890 181116 133962
rect 181076 133884 181128 133890
rect 181076 133826 181128 133832
rect 181168 124228 181220 124234
rect 181168 124170 181220 124176
rect 181180 116006 181208 124170
rect 181168 116000 181220 116006
rect 181168 115942 181220 115948
rect 180984 114572 181036 114578
rect 180984 114514 181036 114520
rect 180996 114442 181024 114514
rect 180984 114436 181036 114442
rect 180984 114378 181036 114384
rect 181168 104916 181220 104922
rect 181168 104858 181220 104864
rect 181180 104802 181208 104858
rect 181088 104774 181208 104802
rect 181088 99414 181116 104774
rect 181076 99408 181128 99414
rect 181076 99350 181128 99356
rect 181168 99340 181220 99346
rect 181168 99282 181220 99288
rect 181180 95282 181208 99282
rect 181088 95254 181208 95282
rect 181088 95198 181116 95254
rect 181076 95192 181128 95198
rect 181076 95134 181128 95140
rect 181168 85604 181220 85610
rect 181168 85546 181220 85552
rect 181180 85490 181208 85546
rect 181088 85462 181208 85490
rect 181088 80102 181116 85462
rect 181076 80096 181128 80102
rect 181076 80038 181128 80044
rect 181168 80028 181220 80034
rect 181168 79970 181220 79976
rect 181180 75970 181208 79970
rect 181088 75942 181208 75970
rect 181088 75886 181116 75942
rect 181076 75880 181128 75886
rect 181076 75822 181128 75828
rect 181168 66292 181220 66298
rect 181168 66234 181220 66240
rect 181180 60858 181208 66234
rect 181168 60852 181220 60858
rect 181168 60794 181220 60800
rect 180984 57928 181036 57934
rect 180984 57870 181036 57876
rect 180996 56574 181024 57870
rect 180984 56568 181036 56574
rect 180984 56510 181036 56516
rect 181168 46980 181220 46986
rect 181168 46922 181220 46928
rect 181180 41478 181208 46922
rect 181168 41472 181220 41478
rect 181168 41414 181220 41420
rect 181076 41404 181128 41410
rect 181076 41346 181128 41352
rect 181088 34746 181116 41346
rect 181076 34740 181128 34746
rect 181076 34682 181128 34688
rect 181168 29028 181220 29034
rect 181168 28970 181220 28976
rect 181180 27606 181208 28970
rect 181168 27600 181220 27606
rect 181168 27542 181220 27548
rect 181168 18012 181220 18018
rect 181168 17954 181220 17960
rect 181180 14550 181208 17954
rect 180984 14544 181036 14550
rect 180984 14486 181036 14492
rect 181168 14544 181220 14550
rect 181168 14486 181220 14492
rect 180996 7954 181024 14486
rect 180984 7948 181036 7954
rect 180984 7890 181036 7896
rect 181352 5296 181404 5302
rect 181352 5238 181404 5244
rect 180892 4548 180944 4554
rect 180892 4490 180944 4496
rect 180800 3732 180852 3738
rect 180800 3674 180852 3680
rect 181364 480 181392 5238
rect 182192 3670 182220 175086
rect 182560 171068 182588 175086
rect 182284 171040 182588 171068
rect 182284 4486 182312 171040
rect 183204 164286 183232 175086
rect 182456 164280 182508 164286
rect 182456 164222 182508 164228
rect 183192 164280 183244 164286
rect 183192 164222 183244 164228
rect 182468 157434 182496 164222
rect 182468 157406 182588 157434
rect 182560 157298 182588 157406
rect 182468 157270 182588 157298
rect 182468 125594 182496 157270
rect 182364 125588 182416 125594
rect 182364 125530 182416 125536
rect 182456 125588 182508 125594
rect 182456 125530 182508 125536
rect 182376 114458 182404 125530
rect 182376 114430 182496 114458
rect 182468 104922 182496 114430
rect 182456 104916 182508 104922
rect 182456 104858 182508 104864
rect 182364 103624 182416 103630
rect 182416 103572 182496 103578
rect 182364 103566 182496 103572
rect 182376 103550 182496 103566
rect 182468 102134 182496 103550
rect 182456 102128 182508 102134
rect 182456 102070 182508 102076
rect 182456 97300 182508 97306
rect 182456 97242 182508 97248
rect 182468 84182 182496 97242
rect 182456 84176 182508 84182
rect 182456 84118 182508 84124
rect 182456 79348 182508 79354
rect 182456 79290 182508 79296
rect 182468 66298 182496 79290
rect 182364 66292 182416 66298
rect 182364 66234 182416 66240
rect 182456 66292 182508 66298
rect 182456 66234 182508 66240
rect 182376 64870 182404 66234
rect 182364 64864 182416 64870
rect 182364 64806 182416 64812
rect 182364 48340 182416 48346
rect 182364 48282 182416 48288
rect 182376 46918 182404 48282
rect 182364 46912 182416 46918
rect 182364 46854 182416 46860
rect 182364 37324 182416 37330
rect 182364 37266 182416 37272
rect 182376 31754 182404 37266
rect 182364 31748 182416 31754
rect 182364 31690 182416 31696
rect 182364 29028 182416 29034
rect 182364 28970 182416 28976
rect 182376 22166 182404 28970
rect 183468 28280 183520 28286
rect 183468 28222 183520 28228
rect 182364 22160 182416 22166
rect 182364 22102 182416 22108
rect 182456 22024 182508 22030
rect 182456 21966 182508 21972
rect 182468 14498 182496 21966
rect 182376 14470 182496 14498
rect 182376 8022 182404 14470
rect 182364 8016 182416 8022
rect 182364 7958 182416 7964
rect 182272 4480 182324 4486
rect 182272 4422 182324 4428
rect 183480 4010 183508 28222
rect 182548 4004 182600 4010
rect 182548 3946 182600 3952
rect 183468 4004 183520 4010
rect 183468 3946 183520 3952
rect 182180 3664 182232 3670
rect 182180 3606 182232 3612
rect 182560 480 182588 3946
rect 183572 3806 183600 175086
rect 184032 171068 184060 175086
rect 183664 171040 184060 171068
rect 183664 4418 183692 171040
rect 184492 164286 184520 175222
rect 184952 175086 185334 175114
rect 183928 164280 183980 164286
rect 183928 164222 183980 164228
rect 184480 164280 184532 164286
rect 184480 164222 184532 164228
rect 183940 153406 183968 164222
rect 183928 153400 183980 153406
rect 183928 153342 183980 153348
rect 183928 153264 183980 153270
rect 183928 153206 183980 153212
rect 183940 143546 183968 153206
rect 183928 143540 183980 143546
rect 183928 143482 183980 143488
rect 183928 124296 183980 124302
rect 183848 124244 183928 124250
rect 183848 124238 183980 124244
rect 183848 124222 183968 124238
rect 183848 122806 183876 124222
rect 183836 122800 183888 122806
rect 183836 122742 183888 122748
rect 183928 113212 183980 113218
rect 183928 113154 183980 113160
rect 183940 104922 183968 113154
rect 183836 104916 183888 104922
rect 183836 104858 183888 104864
rect 183928 104916 183980 104922
rect 183928 104858 183980 104864
rect 183848 101454 183876 104858
rect 183836 101448 183888 101454
rect 183836 101390 183888 101396
rect 183836 101312 183888 101318
rect 183836 101254 183888 101260
rect 183848 85814 183876 101254
rect 183836 85808 183888 85814
rect 183836 85750 183888 85756
rect 183836 84244 183888 84250
rect 183836 84186 183888 84192
rect 183848 84130 183876 84186
rect 183848 84102 183968 84130
rect 183940 74769 183968 84102
rect 183926 74760 183982 74769
rect 183926 74695 183982 74704
rect 183834 74624 183890 74633
rect 183834 74559 183890 74568
rect 183848 70718 183876 74559
rect 183836 70712 183888 70718
rect 183836 70654 183888 70660
rect 183836 66292 183888 66298
rect 183836 66234 183888 66240
rect 183848 64870 183876 66234
rect 183836 64864 183888 64870
rect 183836 64806 183888 64812
rect 183836 55276 183888 55282
rect 183836 55218 183888 55224
rect 183848 50402 183876 55218
rect 183848 50374 183968 50402
rect 183940 45626 183968 50374
rect 183928 45620 183980 45626
rect 183928 45562 183980 45568
rect 184020 45620 184072 45626
rect 184020 45562 184072 45568
rect 184032 35986 184060 45562
rect 183940 35958 184060 35986
rect 183940 27742 183968 35958
rect 183928 27736 183980 27742
rect 183928 27678 183980 27684
rect 183744 26376 183796 26382
rect 183744 26318 183796 26324
rect 183756 26246 183784 26318
rect 183744 26240 183796 26246
rect 183744 26182 183796 26188
rect 183744 16652 183796 16658
rect 183744 16594 183796 16600
rect 183756 13190 183784 16594
rect 184848 14476 184900 14482
rect 184848 14418 184900 14424
rect 183744 13184 183796 13190
rect 183744 13126 183796 13132
rect 184756 9036 184808 9042
rect 184756 8978 184808 8984
rect 183652 4412 183704 4418
rect 183652 4354 183704 4360
rect 183560 3800 183612 3806
rect 183560 3742 183612 3748
rect 183744 3528 183796 3534
rect 183744 3470 183796 3476
rect 183756 480 183784 3470
rect 184768 3346 184796 8978
rect 184860 3534 184888 14418
rect 184952 3874 184980 175086
rect 185412 172514 185440 175222
rect 186346 175086 186544 175114
rect 185124 172508 185176 172514
rect 185124 172450 185176 172456
rect 185400 172508 185452 172514
rect 185400 172450 185452 172456
rect 185136 162897 185164 172450
rect 186412 171080 186464 171086
rect 186412 171022 186464 171028
rect 186320 171012 186372 171018
rect 186320 170954 186372 170960
rect 185122 162888 185178 162897
rect 185122 162823 185178 162832
rect 185306 162888 185362 162897
rect 185306 162823 185362 162832
rect 185320 153270 185348 162823
rect 185216 153264 185268 153270
rect 185216 153206 185268 153212
rect 185308 153264 185360 153270
rect 185308 153206 185360 153212
rect 185228 148458 185256 153206
rect 185228 148430 185440 148458
rect 185412 137850 185440 148430
rect 185228 137822 185440 137850
rect 185228 116006 185256 137822
rect 185124 116000 185176 116006
rect 185124 115942 185176 115948
rect 185216 116000 185268 116006
rect 185216 115942 185268 115948
rect 185136 114510 185164 115942
rect 185124 114504 185176 114510
rect 185124 114446 185176 114452
rect 185216 111036 185268 111042
rect 185216 110978 185268 110984
rect 185228 96626 185256 110978
rect 185032 96620 185084 96626
rect 185032 96562 185084 96568
rect 185216 96620 185268 96626
rect 185216 96562 185268 96568
rect 185044 95198 185072 96562
rect 185032 95192 185084 95198
rect 185032 95134 185084 95140
rect 185216 85604 185268 85610
rect 185216 85546 185268 85552
rect 185228 77330 185256 85546
rect 185136 77302 185256 77330
rect 185136 70446 185164 77302
rect 185124 70440 185176 70446
rect 185124 70382 185176 70388
rect 185216 70304 185268 70310
rect 185216 70246 185268 70252
rect 185228 64870 185256 70246
rect 185216 64864 185268 64870
rect 185216 64806 185268 64812
rect 185124 59220 185176 59226
rect 185124 59162 185176 59168
rect 185136 45558 185164 59162
rect 185124 45552 185176 45558
rect 185124 45494 185176 45500
rect 185400 45552 185452 45558
rect 185400 45494 185452 45500
rect 185412 18018 185440 45494
rect 186228 26920 186280 26926
rect 186228 26862 186280 26868
rect 185124 18012 185176 18018
rect 185124 17954 185176 17960
rect 185400 18012 185452 18018
rect 185400 17954 185452 17960
rect 185136 12510 185164 17954
rect 185124 12504 185176 12510
rect 185124 12446 185176 12452
rect 184940 3868 184992 3874
rect 184940 3810 184992 3816
rect 184848 3528 184900 3534
rect 184848 3470 184900 3476
rect 184768 3318 184888 3346
rect 184860 480 184888 3318
rect 186240 626 186268 26862
rect 186332 4078 186360 170954
rect 186424 4282 186452 171022
rect 186516 8158 186544 175086
rect 186608 175086 186806 175114
rect 186976 175086 187266 175114
rect 187818 175086 188108 175114
rect 186608 171018 186636 175086
rect 186976 171086 187004 175086
rect 188080 174010 188108 175086
rect 188172 175086 188278 175114
rect 188448 175086 188738 175114
rect 189198 175086 189304 175114
rect 188068 174004 188120 174010
rect 188068 173946 188120 173952
rect 186964 171080 187016 171086
rect 186964 171022 187016 171028
rect 187792 171080 187844 171086
rect 187792 171022 187844 171028
rect 186596 171012 186648 171018
rect 186596 170954 186648 170960
rect 187700 169448 187752 169454
rect 187700 169390 187752 169396
rect 187608 15904 187660 15910
rect 187608 15846 187660 15852
rect 186504 8152 186556 8158
rect 186504 8094 186556 8100
rect 186412 4276 186464 4282
rect 186412 4218 186464 4224
rect 186320 4072 186372 4078
rect 186320 4014 186372 4020
rect 186056 598 186268 626
rect 187620 610 187648 15846
rect 187712 4146 187740 169390
rect 187804 6594 187832 171022
rect 188172 169454 188200 175086
rect 188448 171086 188476 175086
rect 188436 171080 188488 171086
rect 188436 171022 188488 171028
rect 189080 171080 189132 171086
rect 189080 171022 189132 171028
rect 188160 169448 188212 169454
rect 188160 169390 188212 169396
rect 188160 169312 188212 169318
rect 188160 169254 188212 169260
rect 188172 157434 188200 169254
rect 188172 157406 188292 157434
rect 188264 153882 188292 157406
rect 188252 153876 188304 153882
rect 188252 153818 188304 153824
rect 188988 21412 189040 21418
rect 188988 21354 189040 21360
rect 187792 6588 187844 6594
rect 187792 6530 187844 6536
rect 189000 4146 189028 21354
rect 187700 4140 187752 4146
rect 187700 4082 187752 4088
rect 188436 4140 188488 4146
rect 188436 4082 188488 4088
rect 188988 4140 189040 4146
rect 188988 4082 189040 4088
rect 187240 604 187292 610
rect 186056 480 186084 598
rect 187240 546 187292 552
rect 187608 604 187660 610
rect 187608 546 187660 552
rect 187252 480 187280 546
rect 188448 480 188476 4082
rect 189092 3398 189120 171022
rect 189172 171012 189224 171018
rect 189172 170954 189224 170960
rect 189184 6662 189212 170954
rect 189276 152522 189304 175086
rect 189368 175086 189658 175114
rect 189920 175086 190210 175114
rect 189368 171086 189396 175086
rect 189356 171080 189408 171086
rect 189356 171022 189408 171028
rect 189920 171018 189948 175086
rect 190552 171080 190604 171086
rect 190552 171022 190604 171028
rect 189908 171012 189960 171018
rect 189908 170954 189960 170960
rect 189264 152516 189316 152522
rect 189264 152458 189316 152464
rect 190564 6730 190592 171022
rect 190656 151094 190684 175100
rect 190748 175086 191130 175114
rect 191208 175086 191590 175114
rect 190644 151088 190696 151094
rect 190644 151030 190696 151036
rect 190552 6724 190604 6730
rect 190552 6666 190604 6672
rect 189172 6656 189224 6662
rect 189172 6598 189224 6604
rect 189632 3460 189684 3466
rect 189632 3402 189684 3408
rect 189080 3392 189132 3398
rect 189080 3334 189132 3340
rect 189644 480 189672 3402
rect 190748 3330 190776 175086
rect 191208 171086 191236 175086
rect 191196 171080 191248 171086
rect 191196 171022 191248 171028
rect 191932 171080 191984 171086
rect 191932 171022 191984 171028
rect 191944 8226 191972 171022
rect 192036 149734 192064 175100
rect 192128 175086 192602 175114
rect 192680 175086 193062 175114
rect 192024 149728 192076 149734
rect 192024 149670 192076 149676
rect 192024 10396 192076 10402
rect 192024 10338 192076 10344
rect 191932 8220 191984 8226
rect 191932 8162 191984 8168
rect 190828 5432 190880 5438
rect 190828 5374 190880 5380
rect 190736 3324 190788 3330
rect 190736 3266 190788 3272
rect 190840 480 190868 5374
rect 192036 480 192064 10338
rect 192128 3262 192156 175086
rect 192680 171086 192708 175086
rect 193402 173904 193458 173913
rect 193402 173839 193458 173848
rect 192668 171080 192720 171086
rect 192668 171022 192720 171028
rect 193312 171080 193364 171086
rect 193312 171022 193364 171028
rect 193324 7546 193352 171022
rect 193416 164257 193444 173839
rect 193508 169046 193536 175100
rect 193692 175086 193982 175114
rect 194152 175086 194442 175114
rect 194796 175086 194994 175114
rect 195072 175086 195454 175114
rect 195624 175086 195914 175114
rect 196084 175086 196374 175114
rect 193692 173913 193720 175086
rect 193678 173904 193734 173913
rect 193678 173839 193734 173848
rect 194152 171086 194180 175086
rect 194416 173188 194468 173194
rect 194416 173130 194468 173136
rect 194140 171080 194192 171086
rect 194140 171022 194192 171028
rect 193496 169040 193548 169046
rect 193496 168982 193548 168988
rect 193402 164248 193458 164257
rect 193402 164183 193458 164192
rect 193586 164248 193642 164257
rect 193586 164183 193642 164192
rect 193600 154737 193628 164183
rect 193586 154728 193642 154737
rect 193586 154663 193642 154672
rect 193494 154592 193550 154601
rect 193494 154527 193550 154536
rect 193508 144906 193536 154527
rect 193496 144900 193548 144906
rect 193496 144842 193548 144848
rect 193588 144900 193640 144906
rect 193588 144842 193640 144848
rect 193600 128382 193628 144842
rect 194138 144800 194194 144809
rect 194138 144735 194194 144744
rect 194152 144226 194180 144735
rect 194140 144220 194192 144226
rect 194140 144162 194192 144168
rect 193404 128376 193456 128382
rect 193404 128318 193456 128324
rect 193588 128376 193640 128382
rect 193588 128318 193640 128324
rect 193416 118674 193444 128318
rect 193416 118646 193628 118674
rect 193600 109070 193628 118646
rect 193404 109064 193456 109070
rect 193404 109006 193456 109012
rect 193588 109064 193640 109070
rect 193588 109006 193640 109012
rect 193416 99362 193444 109006
rect 193416 99334 193628 99362
rect 193600 89758 193628 99334
rect 193404 89752 193456 89758
rect 193404 89694 193456 89700
rect 193588 89752 193640 89758
rect 193588 89694 193640 89700
rect 193416 80050 193444 89694
rect 193416 80022 193628 80050
rect 193600 57934 193628 80022
rect 193588 57928 193640 57934
rect 193588 57870 193640 57876
rect 193496 48340 193548 48346
rect 193496 48282 193548 48288
rect 193508 41426 193536 48282
rect 193508 41398 193628 41426
rect 193600 31770 193628 41398
rect 193416 31742 193628 31770
rect 193312 7540 193364 7546
rect 193312 7482 193364 7488
rect 193220 3664 193272 3670
rect 193220 3606 193272 3612
rect 192116 3256 192168 3262
rect 192116 3198 192168 3204
rect 193232 480 193260 3606
rect 193416 3194 193444 31742
rect 194428 3670 194456 173130
rect 194692 171080 194744 171086
rect 194692 171022 194744 171028
rect 194600 167884 194652 167890
rect 194600 167826 194652 167832
rect 194508 5364 194560 5370
rect 194508 5306 194560 5312
rect 194416 3664 194468 3670
rect 194416 3606 194468 3612
rect 193404 3188 193456 3194
rect 193404 3130 193456 3136
rect 194520 2666 194548 5306
rect 194612 3126 194640 167826
rect 194704 7478 194732 171022
rect 194796 148374 194824 175086
rect 195072 167890 195100 175086
rect 195624 171086 195652 175086
rect 195612 171080 195664 171086
rect 195612 171022 195664 171028
rect 195060 167884 195112 167890
rect 195060 167826 195112 167832
rect 194784 148368 194836 148374
rect 194784 148310 194836 148316
rect 196084 146946 196112 175086
rect 196452 171068 196480 175222
rect 197386 175086 197492 175114
rect 197268 173256 197320 173262
rect 197268 173198 197320 173204
rect 196176 171040 196480 171068
rect 196176 159066 196204 171040
rect 196176 159038 196296 159066
rect 196072 146940 196124 146946
rect 196072 146882 196124 146888
rect 196268 135425 196296 159038
rect 196254 135416 196310 135425
rect 196254 135351 196310 135360
rect 196162 135280 196218 135289
rect 196162 135215 196218 135224
rect 196176 125594 196204 135215
rect 196164 125588 196216 125594
rect 196164 125530 196216 125536
rect 196164 116000 196216 116006
rect 196164 115942 196216 115948
rect 196176 106282 196204 115942
rect 196164 106276 196216 106282
rect 196164 106218 196216 106224
rect 196164 96688 196216 96694
rect 196164 96630 196216 96636
rect 194692 7472 194744 7478
rect 194692 7414 194744 7420
rect 194600 3120 194652 3126
rect 194600 3062 194652 3068
rect 196176 3058 196204 96630
rect 197280 3058 197308 173198
rect 197464 7410 197492 175086
rect 197556 175086 197846 175114
rect 197556 145586 197584 175086
rect 197924 171068 197952 175222
rect 198766 175086 198964 175114
rect 197648 171040 197952 171068
rect 197648 159066 197676 171040
rect 197648 159038 197768 159066
rect 197544 145580 197596 145586
rect 197544 145522 197596 145528
rect 197740 138122 197768 159038
rect 198936 157554 198964 175086
rect 199028 175086 199226 175114
rect 198924 157548 198976 157554
rect 198924 157490 198976 157496
rect 198924 157344 198976 157350
rect 198924 157286 198976 157292
rect 198738 154592 198794 154601
rect 198738 154527 198794 154536
rect 198752 145081 198780 154527
rect 198738 145072 198794 145081
rect 198738 145007 198794 145016
rect 197740 138094 197860 138122
rect 197832 135289 197860 138094
rect 197634 135280 197690 135289
rect 197634 135215 197690 135224
rect 197818 135280 197874 135289
rect 197818 135215 197874 135224
rect 197648 125594 197676 135215
rect 197636 125588 197688 125594
rect 197636 125530 197688 125536
rect 197636 116000 197688 116006
rect 197636 115942 197688 115948
rect 197648 106282 197676 115942
rect 197636 106276 197688 106282
rect 197636 106218 197688 106224
rect 197636 96688 197688 96694
rect 197636 96630 197688 96636
rect 197452 7404 197504 7410
rect 197452 7346 197504 7352
rect 196164 3052 196216 3058
rect 196164 2994 196216 3000
rect 196808 3052 196860 3058
rect 196808 2994 196860 3000
rect 197268 3052 197320 3058
rect 197268 2994 197320 3000
rect 194428 2638 194548 2666
rect 194428 480 194456 2638
rect 195612 1896 195664 1902
rect 195612 1838 195664 1844
rect 195624 480 195652 1838
rect 196820 480 196848 2994
rect 197648 2990 197676 96630
rect 198936 7342 198964 157286
rect 199028 154601 199056 175086
rect 199764 173602 199792 175100
rect 199752 173596 199804 173602
rect 199752 173538 199804 173544
rect 200028 173324 200080 173330
rect 200028 173266 200080 173272
rect 199014 154592 199070 154601
rect 199014 154527 199070 154536
rect 198924 7336 198976 7342
rect 198924 7278 198976 7284
rect 198004 5500 198056 5506
rect 198004 5442 198056 5448
rect 197636 2984 197688 2990
rect 197636 2926 197688 2932
rect 198016 480 198044 5442
rect 200040 4146 200068 173266
rect 200224 7274 200252 175100
rect 200684 171834 200712 175100
rect 200868 175086 201158 175114
rect 201512 175086 201618 175114
rect 201880 175086 202170 175114
rect 200672 171828 200724 171834
rect 200672 171770 200724 171776
rect 200868 171068 200896 175086
rect 201408 173460 201460 173466
rect 201408 173402 201460 173408
rect 200408 171040 200896 171068
rect 200408 154737 200436 171040
rect 200394 154728 200450 154737
rect 200394 154663 200450 154672
rect 200394 154592 200450 154601
rect 200394 154527 200450 154536
rect 200408 144906 200436 154527
rect 200304 144900 200356 144906
rect 200304 144842 200356 144848
rect 200396 144900 200448 144906
rect 200396 144842 200448 144848
rect 200316 106282 200344 144842
rect 200304 106276 200356 106282
rect 200304 106218 200356 106224
rect 200304 106140 200356 106146
rect 200304 106082 200356 106088
rect 200316 86970 200344 106082
rect 200304 86964 200356 86970
rect 200304 86906 200356 86912
rect 200304 86828 200356 86834
rect 200304 86770 200356 86776
rect 200316 22098 200344 86770
rect 200304 22092 200356 22098
rect 200304 22034 200356 22040
rect 200396 22024 200448 22030
rect 200396 21966 200448 21972
rect 200408 19310 200436 21966
rect 200396 19304 200448 19310
rect 200396 19246 200448 19252
rect 200396 9716 200448 9722
rect 200396 9658 200448 9664
rect 200212 7268 200264 7274
rect 200212 7210 200264 7216
rect 200408 4298 200436 9658
rect 200316 4270 200436 4298
rect 199200 4140 199252 4146
rect 199200 4082 199252 4088
rect 200028 4140 200080 4146
rect 200028 4082 200080 4088
rect 199212 480 199240 4082
rect 200316 2922 200344 4270
rect 201420 4146 201448 173402
rect 201512 167074 201540 175086
rect 201500 167068 201552 167074
rect 201500 167010 201552 167016
rect 201684 167068 201736 167074
rect 201684 167010 201736 167016
rect 201696 162178 201724 167010
rect 201684 162172 201736 162178
rect 201684 162114 201736 162120
rect 201684 161968 201736 161974
rect 201684 161910 201736 161916
rect 201500 159452 201552 159458
rect 201500 159394 201552 159400
rect 201512 142866 201540 159394
rect 201500 142860 201552 142866
rect 201500 142802 201552 142808
rect 201500 7608 201552 7614
rect 201500 7550 201552 7556
rect 200396 4140 200448 4146
rect 200396 4082 200448 4088
rect 201408 4140 201460 4146
rect 201408 4082 201460 4088
rect 200304 2916 200356 2922
rect 200304 2858 200356 2864
rect 200408 480 200436 4082
rect 201512 480 201540 7550
rect 201696 7206 201724 161910
rect 201880 159458 201908 175086
rect 202616 173670 202644 175100
rect 202604 173664 202656 173670
rect 202604 173606 202656 173612
rect 202788 173392 202840 173398
rect 202788 173334 202840 173340
rect 201868 159452 201920 159458
rect 201868 159394 201920 159400
rect 201684 7200 201736 7206
rect 201684 7142 201736 7148
rect 202800 626 202828 173334
rect 202972 171080 203024 171086
rect 202972 171022 203024 171028
rect 202984 141438 203012 171022
rect 202972 141432 203024 141438
rect 202972 141374 203024 141380
rect 203076 7138 203104 175100
rect 203168 175086 203550 175114
rect 203168 171086 203196 175086
rect 204088 173738 204116 175100
rect 204364 175086 204562 175114
rect 204732 175086 205022 175114
rect 205192 175086 205482 175114
rect 204076 173732 204128 173738
rect 204076 173674 204128 173680
rect 204168 173528 204220 173534
rect 204168 173470 204220 173476
rect 203156 171080 203208 171086
rect 203156 171022 203208 171028
rect 203064 7132 203116 7138
rect 203064 7074 203116 7080
rect 204180 626 204208 173470
rect 204260 171080 204312 171086
rect 204260 171022 204312 171028
rect 204272 2854 204300 171022
rect 204364 7070 204392 175086
rect 204732 171068 204760 175086
rect 205192 171086 205220 175086
rect 205928 171902 205956 175100
rect 206020 175086 206494 175114
rect 205916 171896 205968 171902
rect 205916 171838 205968 171844
rect 204548 171040 204760 171068
rect 205180 171080 205232 171086
rect 204548 140078 204576 171040
rect 206020 171034 206048 175086
rect 205180 171022 205232 171028
rect 205744 171006 206048 171034
rect 205744 159390 205772 171006
rect 206572 164257 206600 175222
rect 207032 175086 207414 175114
rect 207492 175086 207874 175114
rect 208044 175086 208334 175114
rect 208504 175086 208886 175114
rect 209056 175086 209346 175114
rect 209806 175086 210188 175114
rect 206928 173596 206980 173602
rect 206928 173538 206980 173544
rect 206006 164248 206062 164257
rect 206006 164183 206008 164192
rect 206060 164183 206062 164192
rect 206558 164248 206614 164257
rect 206558 164183 206614 164192
rect 206008 164154 206060 164160
rect 205732 159384 205784 159390
rect 205732 159326 205784 159332
rect 206008 154624 206060 154630
rect 206008 154566 206060 154572
rect 206020 147694 206048 154566
rect 206008 147688 206060 147694
rect 206008 147630 206060 147636
rect 206100 147620 206152 147626
rect 206100 147562 206152 147568
rect 204536 140072 204588 140078
rect 204536 140014 204588 140020
rect 206112 138038 206140 147562
rect 205916 138032 205968 138038
rect 205916 137974 205968 137980
rect 206100 138032 206152 138038
rect 206100 137974 206152 137980
rect 205928 128382 205956 137974
rect 205732 128376 205784 128382
rect 205916 128376 205968 128382
rect 205784 128324 205864 128330
rect 205732 128318 205864 128324
rect 205916 128318 205968 128324
rect 205744 128302 205864 128318
rect 205836 118726 205864 128302
rect 205824 118720 205876 118726
rect 205824 118662 205876 118668
rect 205916 118652 205968 118658
rect 205916 118594 205968 118600
rect 205928 109070 205956 118594
rect 205732 109064 205784 109070
rect 205916 109064 205968 109070
rect 205784 109012 205864 109018
rect 205732 109006 205864 109012
rect 205916 109006 205968 109012
rect 205744 108990 205864 109006
rect 205836 99414 205864 108990
rect 205824 99408 205876 99414
rect 205824 99350 205876 99356
rect 205916 99340 205968 99346
rect 205916 99282 205968 99288
rect 205928 89758 205956 99282
rect 205732 89752 205784 89758
rect 205916 89752 205968 89758
rect 205784 89700 205864 89706
rect 205732 89694 205864 89700
rect 205916 89694 205968 89700
rect 205744 89678 205864 89694
rect 205836 80102 205864 89678
rect 205824 80096 205876 80102
rect 205824 80038 205876 80044
rect 205916 79960 205968 79966
rect 205916 79902 205968 79908
rect 205928 67726 205956 79902
rect 205916 67720 205968 67726
rect 205916 67662 205968 67668
rect 205824 67652 205876 67658
rect 205824 67594 205876 67600
rect 205836 60738 205864 67594
rect 205836 60710 205956 60738
rect 205928 48414 205956 60710
rect 205916 48408 205968 48414
rect 205916 48350 205968 48356
rect 205824 48340 205876 48346
rect 205824 48282 205876 48288
rect 205836 41426 205864 48282
rect 205836 41398 205956 41426
rect 205928 31754 205956 41398
rect 205732 31748 205784 31754
rect 205732 31690 205784 31696
rect 205916 31748 205968 31754
rect 205916 31690 205968 31696
rect 205744 22794 205772 31690
rect 205744 22766 206048 22794
rect 206020 19258 206048 22766
rect 205928 19230 206048 19258
rect 205928 12442 205956 19230
rect 205732 12436 205784 12442
rect 205732 12378 205784 12384
rect 205916 12436 205968 12442
rect 205916 12378 205968 12384
rect 204352 7064 204404 7070
rect 204352 7006 204404 7012
rect 205744 6798 205772 12378
rect 205732 6792 205784 6798
rect 205732 6734 205784 6740
rect 206940 4146 206968 173538
rect 207032 170474 207060 175086
rect 207492 171034 207520 175086
rect 207124 171006 207520 171034
rect 207020 170468 207072 170474
rect 207020 170410 207072 170416
rect 207124 160818 207152 171006
rect 208044 167414 208072 175086
rect 208400 171080 208452 171086
rect 208400 171022 208452 171028
rect 207204 167408 207256 167414
rect 207204 167350 207256 167356
rect 208032 167408 208084 167414
rect 208032 167350 208084 167356
rect 207112 160812 207164 160818
rect 207112 160754 207164 160760
rect 207216 154737 207244 167350
rect 207202 154728 207258 154737
rect 207202 154663 207258 154672
rect 207202 154592 207258 154601
rect 207202 154527 207204 154536
rect 207256 154527 207258 154536
rect 207480 154556 207532 154562
rect 207204 154498 207256 154504
rect 207480 154498 207532 154504
rect 207492 144922 207520 154498
rect 207308 144894 207520 144922
rect 207308 143546 207336 144894
rect 207296 143540 207348 143546
rect 207296 143482 207348 143488
rect 207296 128308 207348 128314
rect 207296 128250 207348 128256
rect 207308 118726 207336 128250
rect 207296 118720 207348 118726
rect 207296 118662 207348 118668
rect 207388 118652 207440 118658
rect 207388 118594 207440 118600
rect 207400 109018 207428 118594
rect 207308 108990 207428 109018
rect 207308 99414 207336 108990
rect 207296 99408 207348 99414
rect 207296 99350 207348 99356
rect 207388 99340 207440 99346
rect 207388 99282 207440 99288
rect 207400 89706 207428 99282
rect 207216 89678 207428 89706
rect 207216 80170 207244 89678
rect 207204 80164 207256 80170
rect 207204 80106 207256 80112
rect 207112 80028 207164 80034
rect 207112 79970 207164 79976
rect 207124 77246 207152 79970
rect 207112 77240 207164 77246
rect 207112 77182 207164 77188
rect 207204 70372 207256 70378
rect 207204 70314 207256 70320
rect 207216 60722 207244 70314
rect 207204 60716 207256 60722
rect 207204 60658 207256 60664
rect 207388 60716 207440 60722
rect 207388 60658 207440 60664
rect 207400 51134 207428 60658
rect 207388 51128 207440 51134
rect 207388 51070 207440 51076
rect 207296 51060 207348 51066
rect 207296 51002 207348 51008
rect 207308 37505 207336 51002
rect 207294 37496 207350 37505
rect 207294 37431 207350 37440
rect 207386 37360 207442 37369
rect 207386 37295 207442 37304
rect 207400 37262 207428 37295
rect 207388 37256 207440 37262
rect 207388 37198 207440 37204
rect 207388 27668 207440 27674
rect 207388 27610 207440 27616
rect 207400 22166 207428 27610
rect 207388 22160 207440 22166
rect 207388 22102 207440 22108
rect 207204 18012 207256 18018
rect 207204 17954 207256 17960
rect 207216 14498 207244 17954
rect 208412 17270 208440 171022
rect 208504 166394 208532 175086
rect 209056 171086 209084 175086
rect 209044 171080 209096 171086
rect 209044 171022 209096 171028
rect 209872 167476 209924 167482
rect 209872 167418 209924 167424
rect 208492 166388 208544 166394
rect 208492 166330 208544 166336
rect 209884 156738 209912 167418
rect 209872 156732 209924 156738
rect 209872 156674 209924 156680
rect 210160 154630 210188 175086
rect 210252 169114 210280 175100
rect 210344 175086 210726 175114
rect 211278 175086 211384 175114
rect 210240 169108 210292 169114
rect 210240 169050 210292 169056
rect 210344 167482 210372 175086
rect 211068 173868 211120 173874
rect 211068 173810 211120 173816
rect 210332 167476 210384 167482
rect 210332 167418 210384 167424
rect 210056 154624 210108 154630
rect 210056 154566 210108 154572
rect 210148 154624 210200 154630
rect 210148 154566 210200 154572
rect 210068 138122 210096 154566
rect 209976 138094 210096 138122
rect 209976 137986 210004 138094
rect 209976 137958 210188 137986
rect 210160 135250 210188 137958
rect 210148 135244 210200 135250
rect 210148 135186 210200 135192
rect 210056 128308 210108 128314
rect 210056 128250 210108 128256
rect 210068 120714 210096 128250
rect 209884 120686 210096 120714
rect 209884 115977 209912 120686
rect 209870 115968 209926 115977
rect 209870 115903 209926 115912
rect 210146 115968 210202 115977
rect 210146 115903 210202 115912
rect 210160 109018 210188 115903
rect 210068 108990 210188 109018
rect 210068 101402 210096 108990
rect 209884 101374 210096 101402
rect 209884 96665 209912 101374
rect 209870 96656 209926 96665
rect 209870 96591 209926 96600
rect 210146 96656 210202 96665
rect 210146 96591 210202 96600
rect 210160 89706 210188 96591
rect 209976 89678 210188 89706
rect 209976 86970 210004 89678
rect 209964 86964 210016 86970
rect 209964 86906 210016 86912
rect 209872 77308 209924 77314
rect 209872 77250 209924 77256
rect 209884 70258 209912 77250
rect 209884 70230 210004 70258
rect 209976 60722 210004 70230
rect 209964 60716 210016 60722
rect 209964 60658 210016 60664
rect 210148 60716 210200 60722
rect 210148 60658 210200 60664
rect 210160 57934 210188 60658
rect 210148 57928 210200 57934
rect 210148 57870 210200 57876
rect 210056 48340 210108 48346
rect 210056 48282 210108 48288
rect 210068 46918 210096 48282
rect 210056 46912 210108 46918
rect 210056 46854 210108 46860
rect 210148 37324 210200 37330
rect 210148 37266 210200 37272
rect 210160 22250 210188 37266
rect 210068 22222 210188 22250
rect 210068 22114 210096 22222
rect 209976 22086 210096 22114
rect 209976 21978 210004 22086
rect 209976 21950 210096 21978
rect 208400 17264 208452 17270
rect 208400 17206 208452 17212
rect 207216 14470 207336 14498
rect 207308 6866 207336 14470
rect 207296 6860 207348 6866
rect 207296 6802 207348 6808
rect 210068 6118 210096 21950
rect 210056 6112 210108 6118
rect 210056 6054 210108 6060
rect 206284 4140 206336 4146
rect 206284 4082 206336 4088
rect 206928 4140 206980 4146
rect 206928 4082 206980 4088
rect 204260 2848 204312 2854
rect 204260 2790 204312 2796
rect 205088 1284 205140 1290
rect 205088 1226 205140 1232
rect 202708 598 202828 626
rect 203904 598 204208 626
rect 202708 480 202736 598
rect 203904 480 203932 598
rect 205100 480 205128 1226
rect 206296 480 206324 4082
rect 208676 4004 208728 4010
rect 208676 3946 208728 3952
rect 207480 3664 207532 3670
rect 207480 3606 207532 3612
rect 207492 480 207520 3606
rect 208688 480 208716 3946
rect 209872 3868 209924 3874
rect 209872 3810 209924 3816
rect 209884 480 209912 3810
rect 211080 480 211108 173810
rect 211252 171080 211304 171086
rect 211252 171022 211304 171028
rect 211264 22778 211292 171022
rect 211252 22772 211304 22778
rect 211252 22714 211304 22720
rect 211356 6050 211384 175086
rect 211724 167754 211752 175100
rect 211816 175086 212198 175114
rect 212552 175086 212658 175114
rect 212736 175086 213118 175114
rect 213288 175086 213670 175114
rect 213932 175086 214130 175114
rect 214300 175086 214590 175114
rect 214760 175086 215050 175114
rect 215312 175086 215510 175114
rect 215588 175086 216062 175114
rect 211816 171086 211844 175086
rect 211804 171080 211856 171086
rect 211804 171022 211856 171028
rect 211712 167748 211764 167754
rect 211712 167690 211764 167696
rect 211344 6044 211396 6050
rect 211344 5986 211396 5992
rect 212552 5982 212580 175086
rect 212632 167952 212684 167958
rect 212632 167894 212684 167900
rect 212644 158098 212672 167894
rect 212736 164898 212764 175086
rect 213288 167958 213316 175086
rect 213828 173732 213880 173738
rect 213828 173674 213880 173680
rect 213276 167952 213328 167958
rect 213276 167894 213328 167900
rect 212724 164892 212776 164898
rect 212724 164834 212776 164840
rect 212632 158092 212684 158098
rect 212632 158034 212684 158040
rect 212540 5976 212592 5982
rect 212540 5918 212592 5924
rect 212264 3460 212316 3466
rect 212264 3402 212316 3408
rect 212276 480 212304 3402
rect 213840 626 213868 173674
rect 213932 5914 213960 175086
rect 214012 171080 214064 171086
rect 214300 171034 214328 175086
rect 214564 173052 214616 173058
rect 214564 172994 214616 173000
rect 214012 171022 214064 171028
rect 214024 155310 214052 171022
rect 214116 171006 214328 171034
rect 214116 163606 214144 171006
rect 214104 163600 214156 163606
rect 214104 163542 214156 163548
rect 214012 155304 214064 155310
rect 214012 155246 214064 155252
rect 214576 24138 214604 172994
rect 214760 171086 214788 175086
rect 214748 171080 214800 171086
rect 214748 171022 214800 171028
rect 215312 167074 215340 175086
rect 215588 171170 215616 175086
rect 216508 173058 216536 175100
rect 216784 175086 216982 175114
rect 216496 173052 216548 173058
rect 216496 172994 216548 173000
rect 216588 173052 216640 173058
rect 216588 172994 216640 173000
rect 215944 172576 215996 172582
rect 215944 172518 215996 172524
rect 215404 171142 215616 171170
rect 215300 167068 215352 167074
rect 215300 167010 215352 167016
rect 215404 162246 215432 171142
rect 215484 167068 215536 167074
rect 215484 167010 215536 167016
rect 215392 162240 215444 162246
rect 215392 162182 215444 162188
rect 214564 24132 214616 24138
rect 214564 24074 214616 24080
rect 213920 5908 213972 5914
rect 213920 5850 213972 5856
rect 215496 5846 215524 167010
rect 215956 25566 215984 172518
rect 215944 25560 215996 25566
rect 215944 25502 215996 25508
rect 215484 5840 215536 5846
rect 215484 5782 215536 5788
rect 216600 4146 216628 172994
rect 216784 5778 216812 175086
rect 217060 169114 217088 175222
rect 217876 173120 217928 173126
rect 217876 173062 217928 173068
rect 217888 170082 217916 173062
rect 217980 172582 218008 175100
rect 218164 175086 218454 175114
rect 218624 175086 218914 175114
rect 219084 175086 219374 175114
rect 219452 175086 219834 175114
rect 217968 172576 218020 172582
rect 217968 172518 218020 172524
rect 218060 170536 218112 170542
rect 218060 170478 218112 170484
rect 217888 170054 218008 170082
rect 217048 169108 217100 169114
rect 217048 169050 217100 169056
rect 217232 169108 217284 169114
rect 217232 169050 217284 169056
rect 217244 164257 217272 169050
rect 217046 164248 217102 164257
rect 216956 164212 217008 164218
rect 217046 164183 217048 164192
rect 216956 164154 217008 164160
rect 217100 164183 217102 164192
rect 217230 164248 217286 164257
rect 217230 164183 217286 164192
rect 217048 164154 217100 164160
rect 216968 159202 216996 164154
rect 216968 159174 217088 159202
rect 217060 145081 217088 159174
rect 217046 145072 217102 145081
rect 217046 145007 217102 145016
rect 217046 144936 217102 144945
rect 217046 144871 217102 144880
rect 217060 138106 217088 144871
rect 217048 138100 217100 138106
rect 217048 138042 217100 138048
rect 217048 137964 217100 137970
rect 217048 137906 217100 137912
rect 217060 125594 217088 137906
rect 216956 125588 217008 125594
rect 216956 125530 217008 125536
rect 217048 125588 217100 125594
rect 217048 125530 217100 125536
rect 216968 106298 216996 125530
rect 216968 106270 217088 106298
rect 217060 99482 217088 106270
rect 217048 99476 217100 99482
rect 217048 99418 217100 99424
rect 217048 96620 217100 96626
rect 217048 96562 217100 96568
rect 217060 86970 217088 96562
rect 216956 86964 217008 86970
rect 216956 86906 217008 86912
rect 217048 86964 217100 86970
rect 217048 86906 217100 86912
rect 216968 72570 216996 86906
rect 216968 72542 217180 72570
rect 217152 70258 217180 72542
rect 217060 70230 217180 70258
rect 217060 67590 217088 70230
rect 217048 67584 217100 67590
rect 217048 67526 217100 67532
rect 217048 56636 217100 56642
rect 217048 56578 217100 56584
rect 217060 56522 217088 56578
rect 216968 56494 217088 56522
rect 216968 29034 216996 56494
rect 216956 29028 217008 29034
rect 216956 28970 217008 28976
rect 217048 29028 217100 29034
rect 217048 28970 217100 28976
rect 217060 27606 217088 28970
rect 217048 27600 217100 27606
rect 217048 27542 217100 27548
rect 216956 9716 217008 9722
rect 216956 9658 217008 9664
rect 216772 5772 216824 5778
rect 216772 5714 216824 5720
rect 216968 4826 216996 9658
rect 216956 4820 217008 4826
rect 216956 4762 217008 4768
rect 217980 4146 218008 170054
rect 218072 4894 218100 170478
rect 218164 6186 218192 175086
rect 218624 170542 218652 175086
rect 218612 170536 218664 170542
rect 218612 170478 218664 170484
rect 219084 170354 219112 175086
rect 219348 173800 219400 173806
rect 219348 173742 219400 173748
rect 218348 170326 219112 170354
rect 218348 154578 218376 170326
rect 218256 154562 218376 154578
rect 218244 154556 218376 154562
rect 218296 154550 218376 154556
rect 218428 154556 218480 154562
rect 218244 154498 218296 154504
rect 218428 154498 218480 154504
rect 218256 154467 218284 154498
rect 218440 149410 218468 154498
rect 218348 149382 218468 149410
rect 218348 130506 218376 149382
rect 218348 130478 218468 130506
rect 218440 125633 218468 130478
rect 218242 125624 218298 125633
rect 218242 125559 218244 125568
rect 218296 125559 218298 125568
rect 218426 125624 218482 125633
rect 218426 125559 218428 125568
rect 218244 125530 218296 125536
rect 218480 125559 218482 125568
rect 218428 125530 218480 125536
rect 218440 119406 218468 125530
rect 218428 119400 218480 119406
rect 218428 119342 218480 119348
rect 218336 114572 218388 114578
rect 218336 114514 218388 114520
rect 218348 106350 218376 114514
rect 218336 106344 218388 106350
rect 218336 106286 218388 106292
rect 218244 106276 218296 106282
rect 218244 106218 218296 106224
rect 218256 104786 218284 106218
rect 218244 104780 218296 104786
rect 218244 104722 218296 104728
rect 218244 100020 218296 100026
rect 218244 99962 218296 99968
rect 218256 95198 218284 99962
rect 218244 95192 218296 95198
rect 218244 95134 218296 95140
rect 218336 91860 218388 91866
rect 218336 91802 218388 91808
rect 218348 75954 218376 91802
rect 218244 75948 218296 75954
rect 218244 75890 218296 75896
rect 218336 75948 218388 75954
rect 218336 75890 218388 75896
rect 218256 66178 218284 75890
rect 218256 66150 218468 66178
rect 218440 56658 218468 66150
rect 218348 56630 218468 56658
rect 218348 56574 218376 56630
rect 218336 56568 218388 56574
rect 218336 56510 218388 56516
rect 218244 46980 218296 46986
rect 218244 46922 218296 46928
rect 218256 38690 218284 46922
rect 218244 38684 218296 38690
rect 218244 38626 218296 38632
rect 218336 38684 218388 38690
rect 218336 38626 218388 38632
rect 218348 29646 218376 38626
rect 218336 29640 218388 29646
rect 218336 29582 218388 29588
rect 218152 6180 218204 6186
rect 218152 6122 218204 6128
rect 218060 4888 218112 4894
rect 218060 4830 218112 4836
rect 215852 4140 215904 4146
rect 215852 4082 215904 4088
rect 216588 4140 216640 4146
rect 216588 4082 216640 4088
rect 217048 4140 217100 4146
rect 217048 4082 217100 4088
rect 217968 4140 218020 4146
rect 217968 4082 218020 4088
rect 218152 4140 218204 4146
rect 218152 4082 218204 4088
rect 214656 3936 214708 3942
rect 214656 3878 214708 3884
rect 213472 598 213868 626
rect 213472 480 213500 598
rect 214668 480 214696 3878
rect 215864 480 215892 4082
rect 217060 480 217088 4082
rect 218164 480 218192 4082
rect 219360 480 219388 173742
rect 219452 6254 219480 175086
rect 219912 171034 219940 175222
rect 219636 171006 219940 171034
rect 219636 154578 219664 171006
rect 219544 154562 219664 154578
rect 219532 154556 219664 154562
rect 219584 154550 219664 154556
rect 219716 154556 219768 154562
rect 219532 154498 219584 154504
rect 219716 154498 219768 154504
rect 219544 154467 219572 154498
rect 219728 149546 219756 154498
rect 219636 149518 219756 149546
rect 219636 143546 219664 149518
rect 219624 143540 219676 143546
rect 219624 143482 219676 143488
rect 219624 134020 219676 134026
rect 219624 133962 219676 133968
rect 219636 133890 219664 133962
rect 219624 133884 219676 133890
rect 219624 133826 219676 133832
rect 219716 133884 219768 133890
rect 219716 133826 219768 133832
rect 219728 119406 219756 133826
rect 219716 119400 219768 119406
rect 219716 119342 219768 119348
rect 219624 114572 219676 114578
rect 219624 114514 219676 114520
rect 219636 104990 219664 114514
rect 219624 104984 219676 104990
rect 219624 104926 219676 104932
rect 219624 104780 219676 104786
rect 219624 104722 219676 104728
rect 219636 98734 219664 104722
rect 219624 98728 219676 98734
rect 219624 98670 219676 98676
rect 219624 75948 219676 75954
rect 219624 75890 219676 75896
rect 219636 72434 219664 75890
rect 219544 72406 219664 72434
rect 219544 58002 219572 72406
rect 219532 57996 219584 58002
rect 219532 57938 219584 57944
rect 219624 57996 219676 58002
rect 219624 57938 219676 57944
rect 219636 48414 219664 57938
rect 219624 48408 219676 48414
rect 219624 48350 219676 48356
rect 219532 48340 219584 48346
rect 219532 48282 219584 48288
rect 219544 38758 219572 48282
rect 219532 38752 219584 38758
rect 219532 38694 219584 38700
rect 219532 35964 219584 35970
rect 219532 35906 219584 35912
rect 219544 27606 219572 35906
rect 219532 27600 219584 27606
rect 219532 27542 219584 27548
rect 219532 9716 219584 9722
rect 219532 9658 219584 9664
rect 219544 8974 219572 9658
rect 219532 8968 219584 8974
rect 219532 8910 219584 8916
rect 219440 6248 219492 6254
rect 219440 6190 219492 6196
rect 220832 4962 220860 175100
rect 220924 175086 221306 175114
rect 221476 175086 221766 175114
rect 220924 5710 220952 175086
rect 221476 173890 221504 175086
rect 221384 173862 221504 173890
rect 221384 162897 221412 173862
rect 221094 162888 221150 162897
rect 221094 162823 221150 162832
rect 221370 162888 221426 162897
rect 221370 162823 221426 162832
rect 221108 130506 221136 162823
rect 221108 130478 221228 130506
rect 221200 125633 221228 130478
rect 221002 125624 221058 125633
rect 221002 125559 221004 125568
rect 221056 125559 221058 125568
rect 221186 125624 221242 125633
rect 221186 125559 221188 125568
rect 221004 125530 221056 125536
rect 221240 125559 221242 125568
rect 221188 125530 221240 125536
rect 221200 117994 221228 125530
rect 221200 117966 221320 117994
rect 221292 113257 221320 117966
rect 221094 113248 221150 113257
rect 221094 113183 221150 113192
rect 221278 113248 221334 113257
rect 221278 113183 221334 113192
rect 221108 106350 221136 113183
rect 221096 106344 221148 106350
rect 221096 106286 221148 106292
rect 221004 106276 221056 106282
rect 221004 106218 221056 106224
rect 221016 85610 221044 106218
rect 221004 85604 221056 85610
rect 221004 85546 221056 85552
rect 221096 85604 221148 85610
rect 221096 85546 221148 85552
rect 221108 66366 221136 85546
rect 221096 66360 221148 66366
rect 221096 66302 221148 66308
rect 221004 66292 221056 66298
rect 221004 66234 221056 66240
rect 221016 58002 221044 66234
rect 221004 57996 221056 58002
rect 221004 57938 221056 57944
rect 221096 57996 221148 58002
rect 221096 57938 221148 57944
rect 221108 48414 221136 57938
rect 221096 48408 221148 48414
rect 221096 48350 221148 48356
rect 221004 48340 221056 48346
rect 221004 48282 221056 48288
rect 221016 46918 221044 48282
rect 221004 46912 221056 46918
rect 221004 46854 221056 46860
rect 221004 37324 221056 37330
rect 221004 37266 221056 37272
rect 221016 27554 221044 37266
rect 221016 27526 221136 27554
rect 221108 22166 221136 27526
rect 221096 22160 221148 22166
rect 221096 22102 221148 22108
rect 221096 22024 221148 22030
rect 221096 21966 221148 21972
rect 221108 10334 221136 21966
rect 221096 10328 221148 10334
rect 221096 10270 221148 10276
rect 220912 5704 220964 5710
rect 220912 5646 220964 5652
rect 222212 5030 222240 175100
rect 222304 175086 222778 175114
rect 222948 175086 223238 175114
rect 223592 175086 223698 175114
rect 223868 175086 224158 175114
rect 222304 5642 222332 175086
rect 222948 164257 222976 175086
rect 223488 172916 223540 172922
rect 223488 172858 223540 172864
rect 222566 164248 222622 164257
rect 222566 164183 222622 164192
rect 222934 164248 222990 164257
rect 222934 164183 222990 164192
rect 222580 133906 222608 164183
rect 222488 133890 222608 133906
rect 222476 133884 222608 133890
rect 222528 133878 222608 133884
rect 222476 133826 222528 133832
rect 222488 133795 222516 133826
rect 222384 124228 222436 124234
rect 222384 124170 222436 124176
rect 222396 115938 222424 124170
rect 222384 115932 222436 115938
rect 222384 115874 222436 115880
rect 222568 115932 222620 115938
rect 222568 115874 222620 115880
rect 222580 106282 222608 115874
rect 222568 106276 222620 106282
rect 222568 106218 222620 106224
rect 222476 96688 222528 96694
rect 222476 96630 222528 96636
rect 222488 89706 222516 96630
rect 222488 89678 222608 89706
rect 222580 77382 222608 89678
rect 222568 77376 222620 77382
rect 222568 77318 222620 77324
rect 222476 77308 222528 77314
rect 222476 77250 222528 77256
rect 222488 73166 222516 77250
rect 222476 73160 222528 73166
rect 222476 73102 222528 73108
rect 222660 63572 222712 63578
rect 222660 63514 222712 63520
rect 222672 54670 222700 63514
rect 222660 54664 222712 54670
rect 222660 54606 222712 54612
rect 222568 45620 222620 45626
rect 222568 45562 222620 45568
rect 222580 28966 222608 45562
rect 222384 28960 222436 28966
rect 222384 28902 222436 28908
rect 222568 28960 222620 28966
rect 222568 28902 222620 28908
rect 222396 19394 222424 28902
rect 222396 19366 222516 19394
rect 222488 19310 222516 19366
rect 222476 19304 222528 19310
rect 222476 19246 222528 19252
rect 222292 5636 222344 5642
rect 222292 5578 222344 5584
rect 222200 5024 222252 5030
rect 222200 4966 222252 4972
rect 220820 4956 220872 4962
rect 220820 4898 220872 4904
rect 223500 4146 223528 172858
rect 223592 5098 223620 175086
rect 223868 171170 223896 175086
rect 224236 172514 224264 175222
rect 224972 175086 225170 175114
rect 225248 175086 225630 175114
rect 224224 172508 224276 172514
rect 224224 172450 224276 172456
rect 223684 171142 223896 171170
rect 223684 6322 223712 171142
rect 223856 162920 223908 162926
rect 223856 162862 223908 162868
rect 223868 157400 223896 162862
rect 223868 157372 223988 157400
rect 223960 151858 223988 157372
rect 223776 151830 223988 151858
rect 223776 151774 223804 151830
rect 223764 151768 223816 151774
rect 223764 151710 223816 151716
rect 223856 142180 223908 142186
rect 223856 142122 223908 142128
rect 223868 124302 223896 142122
rect 223856 124296 223908 124302
rect 223856 124238 223908 124244
rect 223764 122868 223816 122874
rect 223764 122810 223816 122816
rect 223776 116006 223804 122810
rect 223764 116000 223816 116006
rect 223764 115942 223816 115948
rect 223856 115864 223908 115870
rect 223856 115806 223908 115812
rect 223868 103562 223896 115806
rect 223856 103556 223908 103562
rect 223856 103498 223908 103504
rect 223948 103420 224000 103426
rect 223948 103362 224000 103368
rect 223960 85610 223988 103362
rect 223856 85604 223908 85610
rect 223856 85546 223908 85552
rect 223948 85604 224000 85610
rect 223948 85546 224000 85552
rect 223868 64938 223896 85546
rect 223764 64932 223816 64938
rect 223764 64874 223816 64880
rect 223856 64932 223908 64938
rect 223856 64874 223908 64880
rect 223776 58070 223804 64874
rect 223764 58064 223816 58070
rect 223764 58006 223816 58012
rect 223764 57928 223816 57934
rect 223764 57870 223816 57876
rect 223776 48278 223804 57870
rect 223764 48272 223816 48278
rect 223764 48214 223816 48220
rect 223948 48272 224000 48278
rect 223948 48214 224000 48220
rect 223960 27742 223988 48214
rect 223948 27736 224000 27742
rect 223948 27678 224000 27684
rect 223856 27668 223908 27674
rect 223856 27610 223908 27616
rect 223868 18630 223896 27610
rect 223856 18624 223908 18630
rect 223856 18566 223908 18572
rect 223672 6316 223724 6322
rect 223672 6258 223724 6264
rect 224972 5166 225000 175086
rect 225248 171034 225276 175086
rect 226076 171154 226104 175100
rect 226352 175086 226550 175114
rect 226628 175086 227010 175114
rect 225512 171148 225564 171154
rect 225512 171090 225564 171096
rect 226064 171148 226116 171154
rect 226064 171090 226116 171096
rect 225064 171006 225276 171034
rect 225064 6390 225092 171006
rect 225524 162874 225552 171090
rect 225432 162846 225552 162874
rect 225432 161430 225460 162846
rect 225420 161424 225472 161430
rect 225420 161366 225472 161372
rect 225328 151836 225380 151842
rect 225328 151778 225380 151784
rect 225340 147914 225368 151778
rect 225340 147886 225460 147914
rect 225432 143585 225460 147886
rect 225234 143576 225290 143585
rect 225234 143511 225290 143520
rect 225418 143576 225474 143585
rect 225418 143511 225474 143520
rect 225248 133906 225276 143511
rect 225248 133878 225368 133906
rect 225340 124250 225368 133878
rect 225248 124222 225368 124250
rect 225248 116006 225276 124222
rect 225236 116000 225288 116006
rect 225236 115942 225288 115948
rect 225328 115864 225380 115870
rect 225328 115806 225380 115812
rect 225340 111246 225368 115806
rect 225328 111240 225380 111246
rect 225328 111182 225380 111188
rect 225236 111172 225288 111178
rect 225236 111114 225288 111120
rect 225248 106162 225276 111114
rect 225248 106134 225368 106162
rect 225340 66366 225368 106134
rect 225328 66360 225380 66366
rect 225328 66302 225380 66308
rect 225236 66292 225288 66298
rect 225236 66234 225288 66240
rect 225248 58002 225276 66234
rect 225236 57996 225288 58002
rect 225236 57938 225288 57944
rect 225328 57996 225380 58002
rect 225328 57938 225380 57944
rect 225340 53122 225368 57938
rect 225248 53094 225368 53122
rect 225248 48278 225276 53094
rect 225236 48272 225288 48278
rect 225236 48214 225288 48220
rect 225420 48272 225472 48278
rect 225420 48214 225472 48220
rect 225432 30394 225460 48214
rect 225144 30388 225196 30394
rect 225144 30330 225196 30336
rect 225420 30388 225472 30394
rect 225420 30330 225472 30336
rect 225156 13122 225184 30330
rect 225144 13116 225196 13122
rect 225144 13058 225196 13064
rect 225052 6384 225104 6390
rect 225052 6326 225104 6332
rect 226352 5234 226380 175086
rect 226628 171034 226656 175086
rect 226444 171006 226656 171034
rect 226444 6458 226472 171006
rect 227088 164257 227116 175222
rect 227732 175086 228022 175114
rect 228284 175086 228482 175114
rect 228560 175086 228942 175114
rect 229112 175086 229402 175114
rect 227628 172984 227680 172990
rect 227628 172926 227680 172932
rect 226706 164248 226762 164257
rect 226706 164183 226762 164192
rect 227074 164248 227130 164257
rect 227074 164183 227130 164192
rect 226720 157418 226748 164183
rect 226524 157412 226576 157418
rect 226524 157354 226576 157360
rect 226708 157412 226760 157418
rect 226708 157354 226760 157360
rect 226536 147694 226564 157354
rect 226524 147688 226576 147694
rect 226524 147630 226576 147636
rect 226616 147620 226668 147626
rect 226616 147562 226668 147568
rect 226628 138666 226656 147562
rect 226628 138638 226748 138666
rect 226720 128330 226748 138638
rect 226628 128302 226748 128330
rect 226628 118726 226656 128302
rect 226616 118720 226668 118726
rect 226616 118662 226668 118668
rect 226708 118652 226760 118658
rect 226708 118594 226760 118600
rect 226720 109018 226748 118594
rect 226628 108990 226748 109018
rect 226628 100586 226656 108990
rect 226628 100558 226748 100586
rect 226720 66366 226748 100558
rect 226708 66360 226760 66366
rect 226708 66302 226760 66308
rect 226616 66292 226668 66298
rect 226616 66234 226668 66240
rect 226628 46918 226656 66234
rect 226616 46912 226668 46918
rect 226616 46854 226668 46860
rect 226708 46912 226760 46918
rect 226708 46854 226760 46860
rect 226720 31770 226748 46854
rect 226628 31742 226748 31770
rect 226628 28966 226656 31742
rect 226616 28960 226668 28966
rect 226616 28902 226668 28908
rect 226432 6452 226484 6458
rect 226432 6394 226484 6400
rect 226340 5228 226392 5234
rect 226340 5170 226392 5176
rect 224960 5160 225012 5166
rect 224960 5102 225012 5108
rect 223580 5092 223632 5098
rect 223580 5034 223632 5040
rect 222936 4140 222988 4146
rect 222936 4082 222988 4088
rect 223488 4140 223540 4146
rect 223488 4082 223540 4088
rect 221740 4072 221792 4078
rect 221740 4014 221792 4020
rect 220544 4004 220596 4010
rect 220544 3946 220596 3952
rect 220556 480 220584 3946
rect 221752 480 221780 4014
rect 222948 480 222976 4082
rect 227640 3942 227668 172926
rect 227732 5302 227760 175086
rect 227812 171080 227864 171086
rect 227812 171022 227864 171028
rect 227824 14482 227852 171022
rect 228284 164257 228312 175086
rect 228560 171086 228588 175086
rect 229008 172848 229060 172854
rect 229008 172790 229060 172796
rect 228548 171080 228600 171086
rect 228548 171022 228600 171028
rect 227994 164248 228050 164257
rect 227994 164183 228050 164192
rect 228270 164248 228326 164257
rect 228270 164183 228326 164192
rect 228008 147642 228036 164183
rect 228008 147614 228220 147642
rect 228192 133906 228220 147614
rect 228100 133878 228220 133906
rect 228100 115938 228128 133878
rect 228088 115932 228140 115938
rect 228088 115874 228140 115880
rect 228088 106344 228140 106350
rect 228088 106286 228140 106292
rect 228100 98682 228128 106286
rect 228008 98654 228128 98682
rect 228008 92478 228036 98654
rect 227996 92472 228048 92478
rect 227996 92414 228048 92420
rect 228088 82884 228140 82890
rect 228088 82826 228140 82832
rect 228100 77994 228128 82826
rect 228088 77988 228140 77994
rect 228088 77930 228140 77936
rect 227996 64932 228048 64938
rect 227996 64874 228048 64880
rect 228008 55162 228036 64874
rect 228008 55134 228128 55162
rect 228100 28286 228128 55134
rect 228088 28280 228140 28286
rect 228088 28222 228140 28228
rect 227812 14476 227864 14482
rect 227812 14418 227864 14424
rect 227720 5296 227772 5302
rect 227720 5238 227772 5244
rect 226524 3936 226576 3942
rect 226524 3878 226576 3884
rect 227628 3936 227680 3942
rect 227628 3878 227680 3884
rect 225328 3392 225380 3398
rect 225328 3334 225380 3340
rect 224132 3188 224184 3194
rect 224132 3130 224184 3136
rect 224144 480 224172 3130
rect 225340 480 225368 3334
rect 226536 480 226564 3878
rect 229020 3330 229048 172790
rect 229112 9042 229140 175086
rect 229192 171080 229244 171086
rect 229480 171034 229508 175222
rect 230032 175086 230414 175114
rect 230676 175086 230874 175114
rect 230952 175086 231334 175114
rect 231504 175086 231794 175114
rect 231964 175086 232346 175114
rect 230032 171086 230060 175086
rect 229192 171022 229244 171028
rect 229204 15910 229232 171022
rect 229296 171006 229508 171034
rect 230020 171080 230072 171086
rect 230020 171022 230072 171028
rect 230480 171080 230532 171086
rect 230480 171022 230532 171028
rect 229296 26926 229324 171006
rect 229284 26920 229336 26926
rect 229284 26862 229336 26868
rect 229192 15904 229244 15910
rect 229192 15846 229244 15852
rect 229100 9036 229152 9042
rect 229100 8978 229152 8984
rect 230492 5846 230520 171022
rect 230572 171012 230624 171018
rect 230572 170954 230624 170960
rect 230480 5840 230532 5846
rect 230480 5782 230532 5788
rect 230584 5438 230612 170954
rect 230676 21418 230704 175086
rect 230952 171086 230980 175086
rect 231124 172712 231176 172718
rect 231124 172654 231176 172660
rect 230940 171080 230992 171086
rect 230940 171022 230992 171028
rect 230664 21412 230716 21418
rect 230664 21354 230716 21360
rect 230572 5432 230624 5438
rect 230572 5374 230624 5380
rect 231136 3738 231164 172654
rect 231504 171018 231532 175086
rect 231492 171012 231544 171018
rect 231492 170954 231544 170960
rect 231964 10402 231992 175086
rect 232792 173194 232820 175100
rect 233266 175086 233372 175114
rect 232780 173188 232832 173194
rect 232780 173130 232832 173136
rect 232504 172780 232556 172786
rect 232504 172722 232556 172728
rect 231952 10396 232004 10402
rect 231952 10338 232004 10344
rect 230112 3732 230164 3738
rect 230112 3674 230164 3680
rect 231124 3732 231176 3738
rect 231124 3674 231176 3680
rect 227720 3324 227772 3330
rect 227720 3266 227772 3272
rect 229008 3324 229060 3330
rect 229008 3266 229060 3272
rect 227732 480 227760 3266
rect 228916 3256 228968 3262
rect 228916 3198 228968 3204
rect 228928 480 228956 3198
rect 230124 480 230152 3674
rect 232516 3346 232544 172722
rect 233344 5370 233372 175086
rect 233436 175086 233726 175114
rect 233332 5364 233384 5370
rect 233332 5306 233384 5312
rect 233436 4826 233464 175086
rect 234264 172922 234292 175100
rect 234252 172916 234304 172922
rect 234252 172858 234304 172864
rect 234528 172916 234580 172922
rect 234528 172858 234580 172864
rect 233424 4820 233476 4826
rect 233424 4762 233476 4768
rect 234540 3738 234568 172858
rect 234724 5506 234752 175100
rect 235184 173602 235212 175100
rect 235172 173596 235224 173602
rect 235172 173538 235224 173544
rect 235264 173460 235316 173466
rect 235264 173402 235316 173408
rect 234712 5500 234764 5506
rect 234712 5442 234764 5448
rect 234804 4140 234856 4146
rect 234804 4082 234856 4088
rect 233700 3732 233752 3738
rect 233700 3674 233752 3680
rect 234528 3732 234580 3738
rect 234528 3674 234580 3680
rect 232424 3318 232544 3346
rect 232424 3194 232452 3318
rect 232504 3256 232556 3262
rect 232504 3198 232556 3204
rect 232412 3188 232464 3194
rect 232412 3130 232464 3136
rect 231308 2984 231360 2990
rect 231308 2926 231360 2932
rect 231320 480 231348 2926
rect 232516 480 232544 3198
rect 233712 480 233740 3674
rect 234816 480 234844 4082
rect 235276 2990 235304 173402
rect 235644 173398 235672 175100
rect 235632 173392 235684 173398
rect 235632 173334 235684 173340
rect 235908 173324 235960 173330
rect 235908 173266 235960 173272
rect 235920 4146 235948 173266
rect 236104 7614 236132 175100
rect 236656 172650 236684 175100
rect 237116 173262 237144 175100
rect 237104 173256 237156 173262
rect 237104 173198 237156 173204
rect 237288 173256 237340 173262
rect 237288 173198 237340 173204
rect 236644 172644 236696 172650
rect 236644 172586 236696 172592
rect 237300 67946 237328 173198
rect 237472 171080 237524 171086
rect 237472 171022 237524 171028
rect 237208 67918 237328 67946
rect 237208 67674 237236 67918
rect 237208 67646 237328 67674
rect 237300 66230 237328 67646
rect 237288 66224 237340 66230
rect 237288 66166 237340 66172
rect 237288 56636 237340 56642
rect 237288 56578 237340 56584
rect 237300 48634 237328 56578
rect 237208 48606 237328 48634
rect 237208 48346 237236 48606
rect 237196 48340 237248 48346
rect 237196 48282 237248 48288
rect 237288 48340 237340 48346
rect 237288 48282 237340 48288
rect 237300 46918 237328 48282
rect 237288 46912 237340 46918
rect 237288 46854 237340 46860
rect 237288 37324 237340 37330
rect 237288 37266 237340 37272
rect 237300 27606 237328 37266
rect 237288 27600 237340 27606
rect 237288 27542 237340 27548
rect 237196 9716 237248 9722
rect 237196 9658 237248 9664
rect 236092 7608 236144 7614
rect 236092 7550 236144 7556
rect 235908 4140 235960 4146
rect 235908 4082 235960 4088
rect 236000 3256 236052 3262
rect 236000 3198 236052 3204
rect 235264 2984 235316 2990
rect 235264 2926 235316 2932
rect 236012 480 236040 3198
rect 237208 480 237236 9658
rect 237484 3670 237512 171022
rect 237472 3664 237524 3670
rect 237472 3606 237524 3612
rect 237576 3534 237604 175100
rect 238036 172582 238064 175100
rect 238128 175086 238510 175114
rect 238864 175086 239062 175114
rect 239324 175086 239522 175114
rect 238024 172576 238076 172582
rect 238024 172518 238076 172524
rect 238128 171086 238156 175086
rect 238668 173392 238720 173398
rect 238668 173334 238720 173340
rect 238116 171080 238168 171086
rect 238116 171022 238168 171028
rect 238680 67810 238708 173334
rect 238760 122800 238812 122806
rect 238760 122742 238812 122748
rect 238772 106282 238800 122742
rect 238760 106276 238812 106282
rect 238760 106218 238812 106224
rect 238680 67782 238800 67810
rect 238772 67674 238800 67782
rect 238680 67646 238800 67674
rect 238680 66230 238708 67646
rect 238668 66224 238720 66230
rect 238668 66166 238720 66172
rect 238668 56636 238720 56642
rect 238668 56578 238720 56584
rect 238680 48634 238708 56578
rect 238680 48606 238800 48634
rect 238772 48346 238800 48606
rect 238668 48340 238720 48346
rect 238668 48282 238720 48288
rect 238760 48340 238812 48346
rect 238760 48282 238812 48288
rect 238680 46918 238708 48282
rect 238668 46912 238720 46918
rect 238668 46854 238720 46860
rect 238668 37324 238720 37330
rect 238668 37266 238720 37272
rect 238680 27606 238708 37266
rect 238668 27600 238720 27606
rect 238668 27542 238720 27548
rect 238392 9716 238444 9722
rect 238392 9658 238444 9664
rect 237564 3528 237616 3534
rect 237564 3470 237616 3476
rect 238404 480 238432 9658
rect 238864 3806 238892 175086
rect 239324 157434 239352 175086
rect 239968 173670 239996 175100
rect 240244 175086 240442 175114
rect 239956 173664 240008 173670
rect 239956 173606 240008 173612
rect 239048 157406 239352 157434
rect 239048 157298 239076 157406
rect 239048 157270 239168 157298
rect 239140 138122 239168 157270
rect 239048 138094 239168 138122
rect 239048 128382 239076 138094
rect 239036 128376 239088 128382
rect 239036 128318 239088 128324
rect 239128 128308 239180 128314
rect 239128 128250 239180 128256
rect 239140 122806 239168 128250
rect 239128 122800 239180 122806
rect 239128 122742 239180 122748
rect 239036 106276 239088 106282
rect 239036 106218 239088 106224
rect 239048 101454 239076 106218
rect 239036 101448 239088 101454
rect 239036 101390 239088 101396
rect 239036 101312 239088 101318
rect 239036 101254 239088 101260
rect 239048 86970 239076 101254
rect 239036 86964 239088 86970
rect 239036 86906 239088 86912
rect 239036 77308 239088 77314
rect 239036 77250 239088 77256
rect 239048 58290 239076 77250
rect 239048 58262 239168 58290
rect 239140 58018 239168 58262
rect 239048 57990 239168 58018
rect 239048 57934 239076 57990
rect 239036 57928 239088 57934
rect 239036 57870 239088 57876
rect 239036 48340 239088 48346
rect 239036 48282 239088 48288
rect 239048 38758 239076 48282
rect 239036 38752 239088 38758
rect 239036 38694 239088 38700
rect 239036 37324 239088 37330
rect 239036 37266 239088 37272
rect 239048 28966 239076 37266
rect 239036 28960 239088 28966
rect 239036 28902 239088 28908
rect 239036 22772 239088 22778
rect 239036 22714 239088 22720
rect 239048 3874 239076 22714
rect 240244 3942 240272 175086
rect 240888 173738 240916 175100
rect 241164 175086 241454 175114
rect 240876 173732 240928 173738
rect 240876 173674 240928 173680
rect 241164 171086 241192 175086
rect 241900 173806 241928 175100
rect 241888 173800 241940 173806
rect 241888 173742 241940 173748
rect 241428 173528 241480 173534
rect 241428 173470 241480 173476
rect 240508 171080 240560 171086
rect 240508 171022 240560 171028
rect 241152 171080 241204 171086
rect 241152 171022 241204 171028
rect 240520 164218 240548 171022
rect 240508 164212 240560 164218
rect 240508 164154 240560 164160
rect 240508 156324 240560 156330
rect 240508 156266 240560 156272
rect 240520 138174 240548 156266
rect 240508 138168 240560 138174
rect 240508 138110 240560 138116
rect 240416 133952 240468 133958
rect 240416 133894 240468 133900
rect 240428 124166 240456 133894
rect 240416 124160 240468 124166
rect 240416 124102 240468 124108
rect 240416 114572 240468 114578
rect 240416 114514 240468 114520
rect 240428 106282 240456 114514
rect 240416 106276 240468 106282
rect 240416 106218 240468 106224
rect 240416 96688 240468 96694
rect 240416 96630 240468 96636
rect 240428 86970 240456 96630
rect 240416 86964 240468 86970
rect 240416 86906 240468 86912
rect 240416 77308 240468 77314
rect 240416 77250 240468 77256
rect 240428 67590 240456 77250
rect 240416 67584 240468 67590
rect 240416 67526 240468 67532
rect 240416 62756 240468 62762
rect 240416 62698 240468 62704
rect 240428 41426 240456 62698
rect 240336 41398 240456 41426
rect 240336 41290 240364 41398
rect 240336 41262 240456 41290
rect 240428 22114 240456 41262
rect 240336 22086 240456 22114
rect 240336 21978 240364 22086
rect 240336 21950 240456 21978
rect 240232 3936 240284 3942
rect 240232 3878 240284 3884
rect 239036 3868 239088 3874
rect 239036 3810 239088 3816
rect 238852 3800 238904 3806
rect 238852 3742 238904 3748
rect 240428 3602 240456 21950
rect 241440 4146 241468 173470
rect 242360 173126 242388 175100
rect 242348 173120 242400 173126
rect 242348 173062 242400 173068
rect 242452 171034 242480 175222
rect 243280 173874 243308 175100
rect 243556 175086 243846 175114
rect 244306 175086 244412 175114
rect 243268 173868 243320 173874
rect 243268 173810 243320 173816
rect 242808 173664 242860 173670
rect 242808 173606 242860 173612
rect 241624 171006 242480 171034
rect 240784 4140 240836 4146
rect 240784 4082 240836 4088
rect 241428 4140 241480 4146
rect 241428 4082 241480 4088
rect 240416 3596 240468 3602
rect 240416 3538 240468 3544
rect 239588 3460 239640 3466
rect 239588 3402 239640 3408
rect 239600 480 239628 3402
rect 240796 480 240824 4082
rect 241624 4010 241652 171006
rect 241612 4004 241664 4010
rect 241612 3946 241664 3952
rect 242820 3534 242848 173606
rect 243556 172718 243584 175086
rect 243084 172712 243136 172718
rect 243084 172654 243136 172660
rect 243544 172712 243596 172718
rect 243544 172654 243596 172660
rect 243096 157434 243124 172654
rect 243544 172576 243596 172582
rect 243544 172518 243596 172524
rect 242912 157406 243124 157434
rect 242912 157298 242940 157406
rect 242912 157270 243032 157298
rect 243004 157162 243032 157270
rect 243004 157134 243124 157162
rect 243096 138106 243124 157134
rect 243084 138100 243136 138106
rect 243084 138042 243136 138048
rect 242992 138032 243044 138038
rect 242992 137974 243044 137980
rect 243004 128466 243032 137974
rect 242912 128438 243032 128466
rect 242912 128330 242940 128438
rect 242912 128302 243032 128330
rect 243004 109154 243032 128302
rect 242912 109126 243032 109154
rect 242912 109018 242940 109126
rect 242912 108990 243032 109018
rect 243004 89842 243032 108990
rect 242912 89814 243032 89842
rect 242912 89706 242940 89814
rect 242912 89678 243032 89706
rect 243004 70394 243032 89678
rect 242912 70366 243032 70394
rect 242912 70258 242940 70366
rect 242912 70230 243032 70258
rect 243004 51082 243032 70230
rect 242912 51054 243032 51082
rect 242912 50946 242940 51054
rect 242912 50918 243032 50946
rect 243004 31770 243032 50918
rect 242912 31742 243032 31770
rect 242912 31634 242940 31742
rect 242912 31606 243032 31634
rect 243004 12458 243032 31606
rect 242912 12430 243032 12458
rect 242912 3738 242940 12430
rect 243176 4072 243228 4078
rect 243176 4014 243228 4020
rect 242900 3732 242952 3738
rect 242900 3674 242952 3680
rect 241980 3528 242032 3534
rect 241980 3470 242032 3476
rect 242808 3528 242860 3534
rect 242808 3470 242860 3476
rect 241992 480 242020 3470
rect 243188 480 243216 4014
rect 243556 3126 243584 172518
rect 244384 4298 244412 175086
rect 244752 173058 244780 175100
rect 244924 173596 244976 173602
rect 244924 173538 244976 173544
rect 244740 173052 244792 173058
rect 244740 172994 244792 173000
rect 244292 4270 244412 4298
rect 244292 4146 244320 4270
rect 244280 4140 244332 4146
rect 244280 4082 244332 4088
rect 244372 4140 244424 4146
rect 244372 4082 244424 4088
rect 243544 3120 243596 3126
rect 243544 3062 243596 3068
rect 244384 480 244412 4082
rect 244936 4078 244964 173538
rect 245212 172786 245240 175100
rect 245686 175086 245792 175114
rect 245568 173732 245620 173738
rect 245568 173674 245620 173680
rect 245200 172780 245252 172786
rect 245200 172722 245252 172728
rect 245580 4146 245608 173674
rect 245568 4140 245620 4146
rect 245568 4082 245620 4088
rect 244924 4072 244976 4078
rect 244924 4014 244976 4020
rect 245764 3398 245792 175086
rect 246224 172990 246252 175100
rect 246304 173868 246356 173874
rect 246304 173810 246356 173816
rect 246212 172984 246264 172990
rect 246212 172926 246264 172932
rect 245752 3392 245804 3398
rect 245752 3334 245804 3340
rect 246316 2922 246344 173810
rect 246684 172854 246712 175100
rect 246948 173800 247000 173806
rect 246948 173742 247000 173748
rect 246672 172848 246724 172854
rect 246672 172790 246724 172796
rect 246960 4842 246988 173742
rect 246776 4814 246988 4842
rect 245568 2916 245620 2922
rect 245568 2858 245620 2864
rect 246304 2916 246356 2922
rect 246304 2858 246356 2864
rect 245580 480 245608 2858
rect 246776 480 246804 4814
rect 247144 3330 247172 175100
rect 247604 172922 247632 175100
rect 248064 173466 248092 175100
rect 248052 173460 248104 173466
rect 248052 173402 248104 173408
rect 248328 173460 248380 173466
rect 248328 173402 248380 173408
rect 247592 172916 247644 172922
rect 247592 172858 247644 172864
rect 248340 4842 248368 173402
rect 248616 172582 248644 175100
rect 249076 173194 249104 175100
rect 249536 173330 249564 175100
rect 249904 175086 250010 175114
rect 249524 173324 249576 173330
rect 249524 173266 249576 173272
rect 249064 173188 249116 173194
rect 249064 173130 249116 173136
rect 249708 173052 249760 173058
rect 249708 172994 249760 173000
rect 248604 172576 248656 172582
rect 248604 172518 248656 172524
rect 247972 4814 248368 4842
rect 247132 3324 247184 3330
rect 247132 3266 247184 3272
rect 247972 480 248000 4814
rect 249720 3534 249748 172994
rect 249156 3528 249208 3534
rect 249156 3470 249208 3476
rect 249708 3528 249760 3534
rect 249708 3470 249760 3476
rect 249168 480 249196 3470
rect 249904 3466 249932 175086
rect 250548 173262 250576 175100
rect 251008 173398 251036 175100
rect 251376 175086 251482 175114
rect 250996 173392 251048 173398
rect 250996 173334 251048 173340
rect 250536 173256 250588 173262
rect 250536 173198 250588 173204
rect 251088 173188 251140 173194
rect 251088 173130 251140 173136
rect 249892 3460 249944 3466
rect 249892 3402 249944 3408
rect 251100 3126 251128 173130
rect 251376 3670 251404 175086
rect 251928 173534 251956 175100
rect 252388 173670 252416 175100
rect 252376 173664 252428 173670
rect 252376 173606 252428 173612
rect 252940 173602 252968 175100
rect 253400 173738 253428 175100
rect 253860 173874 253888 175100
rect 253848 173868 253900 173874
rect 253848 173810 253900 173816
rect 254320 173806 254348 175100
rect 254308 173800 254360 173806
rect 254308 173742 254360 173748
rect 253388 173732 253440 173738
rect 253388 173674 253440 173680
rect 252928 173596 252980 173602
rect 252928 173538 252980 173544
rect 251916 173528 251968 173534
rect 251916 173470 251968 173476
rect 254780 173466 254808 175100
rect 254768 173460 254820 173466
rect 254768 173402 254820 173408
rect 255332 173058 255360 175100
rect 255792 173194 255820 175100
rect 255780 173188 255832 173194
rect 255780 173130 255832 173136
rect 255320 173052 255372 173058
rect 255320 172994 255372 173000
rect 253848 172712 253900 172718
rect 253848 172654 253900 172660
rect 251364 3664 251416 3670
rect 251364 3606 251416 3612
rect 253860 3534 253888 172654
rect 255228 172644 255280 172650
rect 255228 172586 255280 172592
rect 254584 172576 254636 172582
rect 254584 172518 254636 172524
rect 252652 3528 252704 3534
rect 252652 3470 252704 3476
rect 253848 3528 253900 3534
rect 253848 3470 253900 3476
rect 251456 3256 251508 3262
rect 251456 3198 251508 3204
rect 250352 3120 250404 3126
rect 250352 3062 250404 3068
rect 251088 3120 251140 3126
rect 251088 3062 251140 3068
rect 250364 480 250392 3062
rect 251468 480 251496 3198
rect 252664 480 252692 3470
rect 254596 3262 254624 172518
rect 254584 3256 254636 3262
rect 254584 3198 254636 3204
rect 253848 3188 253900 3194
rect 253848 3130 253900 3136
rect 253860 480 253888 3130
rect 255240 2854 255268 172586
rect 256252 172582 256280 175100
rect 256608 172780 256660 172786
rect 256608 172722 256660 172728
rect 256240 172576 256292 172582
rect 256240 172518 256292 172524
rect 256514 57896 256570 57905
rect 256514 57831 256570 57840
rect 256528 48346 256556 57831
rect 256516 48340 256568 48346
rect 256516 48282 256568 48288
rect 256514 38584 256570 38593
rect 256514 38519 256570 38528
rect 256528 29034 256556 38519
rect 256516 29028 256568 29034
rect 256516 28970 256568 28976
rect 256620 2854 256648 172722
rect 256712 172718 256740 175100
rect 256700 172712 256752 172718
rect 256700 172654 256752 172660
rect 256896 167006 256924 175222
rect 257724 172650 257752 175100
rect 258184 172786 258212 175100
rect 258276 175086 258658 175114
rect 258828 175086 259118 175114
rect 259578 175086 259684 175114
rect 258172 172780 258224 172786
rect 258172 172722 258224 172728
rect 258276 172666 258304 175086
rect 257712 172644 257764 172650
rect 257712 172586 257764 172592
rect 258000 172638 258304 172666
rect 256884 167000 256936 167006
rect 256884 166942 256936 166948
rect 257068 167000 257120 167006
rect 257068 166942 257120 166948
rect 257080 164218 257108 166942
rect 256792 164212 256844 164218
rect 256792 164154 256844 164160
rect 257068 164212 257120 164218
rect 257068 164154 257120 164160
rect 256804 154601 256832 164154
rect 256790 154592 256846 154601
rect 256790 154527 256846 154536
rect 256974 154592 257030 154601
rect 256974 154527 256976 154536
rect 257028 154527 257030 154536
rect 257160 154556 257212 154562
rect 256976 154498 257028 154504
rect 257160 154498 257212 154504
rect 257172 144945 257200 154498
rect 256882 144936 256938 144945
rect 256882 144871 256938 144880
rect 257158 144936 257214 144945
rect 257158 144871 257214 144880
rect 256896 138038 256924 144871
rect 256884 138032 256936 138038
rect 256884 137974 256936 137980
rect 256976 137964 257028 137970
rect 256976 137906 257028 137912
rect 256988 135250 257016 137906
rect 256976 135244 257028 135250
rect 256976 135186 257028 135192
rect 257160 135244 257212 135250
rect 257160 135186 257212 135192
rect 257172 125633 257200 135186
rect 256882 125624 256938 125633
rect 256882 125559 256938 125568
rect 257158 125624 257214 125633
rect 257158 125559 257214 125568
rect 256896 118726 256924 125559
rect 256884 118720 256936 118726
rect 256884 118662 256936 118668
rect 256976 118652 257028 118658
rect 256976 118594 257028 118600
rect 256988 115938 257016 118594
rect 256976 115932 257028 115938
rect 256976 115874 257028 115880
rect 257160 115932 257212 115938
rect 257160 115874 257212 115880
rect 257172 106321 257200 115874
rect 256882 106312 256938 106321
rect 256882 106247 256938 106256
rect 257158 106312 257214 106321
rect 257158 106247 257214 106256
rect 256896 97986 256924 106247
rect 256700 97980 256752 97986
rect 256700 97922 256752 97928
rect 256884 97980 256936 97986
rect 256884 97922 256936 97928
rect 256712 89706 256740 97922
rect 256712 89678 256924 89706
rect 256896 80102 256924 89678
rect 256884 80096 256936 80102
rect 256884 80038 256936 80044
rect 256976 79960 257028 79966
rect 256976 79902 257028 79908
rect 256988 77246 257016 79902
rect 256976 77240 257028 77246
rect 256976 77182 257028 77188
rect 256884 67652 256936 67658
rect 256884 67594 256936 67600
rect 256896 60874 256924 67594
rect 256896 60846 257016 60874
rect 256988 58002 257016 60846
rect 256700 57996 256752 58002
rect 256700 57938 256752 57944
rect 256976 57996 257028 58002
rect 256976 57938 257028 57944
rect 256712 57905 256740 57938
rect 256698 57896 256754 57905
rect 256698 57831 256754 57840
rect 256884 48340 256936 48346
rect 256884 48282 256936 48288
rect 256896 48226 256924 48282
rect 256896 48198 257016 48226
rect 256988 38690 257016 48198
rect 256700 38684 256752 38690
rect 256700 38626 256752 38632
rect 256976 38684 257028 38690
rect 256976 38626 257028 38632
rect 256712 38593 256740 38626
rect 256698 38584 256754 38593
rect 256698 38519 256754 38528
rect 256792 29028 256844 29034
rect 256792 28970 256844 28976
rect 256804 22114 256832 28970
rect 256804 22098 256924 22114
rect 256804 22092 256936 22098
rect 256804 22086 256884 22092
rect 256884 22034 256936 22040
rect 257068 22092 257120 22098
rect 257068 22034 257120 22040
rect 257080 19310 257108 22034
rect 257068 19304 257120 19310
rect 257068 19246 257120 19252
rect 257068 12300 257120 12306
rect 257068 12242 257120 12248
rect 257080 3194 257108 12242
rect 258000 4146 258028 172638
rect 258828 171034 258856 175086
rect 258184 171006 258856 171034
rect 258184 4146 258212 171006
rect 257436 4140 257488 4146
rect 257436 4082 257488 4088
rect 257988 4140 258040 4146
rect 257988 4082 258040 4088
rect 258172 4140 258224 4146
rect 258172 4082 258224 4088
rect 258632 4140 258684 4146
rect 258632 4082 258684 4088
rect 257068 3188 257120 3194
rect 257068 3130 257120 3136
rect 255228 2848 255280 2854
rect 255228 2790 255280 2796
rect 256240 2848 256292 2854
rect 256240 2790 256292 2796
rect 256608 2848 256660 2854
rect 256608 2790 256660 2796
rect 255044 604 255096 610
rect 255044 546 255096 552
rect 255056 480 255084 546
rect 256252 480 256280 2790
rect 257448 480 257476 4082
rect 258644 480 258672 4082
rect 259656 610 259684 175086
rect 260116 172582 260144 175100
rect 260590 175086 260788 175114
rect 260104 172576 260156 172582
rect 260104 172518 260156 172524
rect 260760 4078 260788 175086
rect 261036 172582 261064 175100
rect 261496 172650 261524 175100
rect 261956 173126 261984 175100
rect 262508 173262 262536 175100
rect 262496 173256 262548 173262
rect 262496 173198 262548 173204
rect 261944 173120 261996 173126
rect 261944 173062 261996 173068
rect 262968 172650 262996 175100
rect 263442 175086 263548 175114
rect 261484 172644 261536 172650
rect 261484 172586 261536 172592
rect 262864 172644 262916 172650
rect 262864 172586 262916 172592
rect 262956 172644 263008 172650
rect 262956 172586 263008 172592
rect 260932 172576 260984 172582
rect 260932 172518 260984 172524
rect 261024 172576 261076 172582
rect 261024 172518 261076 172524
rect 262128 172576 262180 172582
rect 262128 172518 262180 172524
rect 260748 4072 260800 4078
rect 260748 4014 260800 4020
rect 260944 626 260972 172518
rect 262140 4146 262168 172518
rect 262128 4140 262180 4146
rect 262128 4082 262180 4088
rect 262220 4072 262272 4078
rect 262220 4014 262272 4020
rect 259644 604 259696 610
rect 259644 546 259696 552
rect 259828 604 259880 610
rect 260944 598 261064 626
rect 259828 546 259880 552
rect 259840 480 259868 546
rect 261036 480 261064 598
rect 262232 480 262260 4014
rect 262876 3058 262904 172586
rect 263416 4140 263468 4146
rect 263416 4082 263468 4088
rect 262864 3052 262916 3058
rect 262864 2994 262916 3000
rect 263428 480 263456 4082
rect 263520 2990 263548 175086
rect 263888 173194 263916 175100
rect 264362 175086 264836 175114
rect 263876 173188 263928 173194
rect 263876 173130 263928 173136
rect 264244 172644 264296 172650
rect 264244 172586 264296 172592
rect 264256 3942 264284 172586
rect 264244 3936 264296 3942
rect 264244 3878 264296 3884
rect 264808 3806 264836 175086
rect 264796 3800 264848 3806
rect 264796 3742 264848 3748
rect 264900 3738 264928 175100
rect 265256 173120 265308 173126
rect 265256 173062 265308 173068
rect 264888 3732 264940 3738
rect 264888 3674 264940 3680
rect 264612 3052 264664 3058
rect 264612 2994 264664 3000
rect 263508 2984 263560 2990
rect 263508 2926 263560 2932
rect 264624 480 264652 2994
rect 265268 610 265296 173062
rect 265360 172786 265388 175100
rect 265348 172780 265400 172786
rect 265348 172722 265400 172728
rect 265820 172650 265848 175100
rect 266176 172780 266228 172786
rect 266176 172722 266228 172728
rect 265808 172644 265860 172650
rect 265808 172586 265860 172592
rect 266188 3670 266216 172722
rect 266176 3664 266228 3670
rect 266176 3606 266228 3612
rect 266280 3602 266308 175100
rect 266544 173256 266596 173262
rect 266544 173198 266596 173204
rect 266268 3596 266320 3602
rect 266268 3538 266320 3544
rect 266556 3346 266584 173198
rect 266832 172786 266860 175100
rect 267306 175086 267596 175114
rect 267004 173188 267056 173194
rect 267004 173130 267056 173136
rect 266820 172780 266872 172786
rect 266820 172722 266872 172728
rect 267016 4010 267044 173130
rect 267004 4004 267056 4010
rect 267004 3946 267056 3952
rect 267568 3466 267596 175086
rect 267752 173126 267780 175100
rect 267740 173120 267792 173126
rect 267740 173062 267792 173068
rect 268212 172786 268240 175100
rect 268686 175086 268884 175114
rect 267648 172780 267700 172786
rect 267648 172722 267700 172728
rect 268200 172780 268252 172786
rect 268200 172722 268252 172728
rect 267660 3534 267688 172722
rect 268384 172644 268436 172650
rect 268384 172586 268436 172592
rect 268108 3936 268160 3942
rect 268108 3878 268160 3884
rect 267648 3528 267700 3534
rect 267648 3470 267700 3476
rect 267556 3460 267608 3466
rect 267556 3402 267608 3408
rect 266556 3318 267044 3346
rect 265256 604 265308 610
rect 265256 546 265308 552
rect 265808 604 265860 610
rect 265808 546 265860 552
rect 265820 480 265848 546
rect 267016 480 267044 3318
rect 268120 480 268148 3878
rect 268396 3330 268424 172586
rect 268856 3874 268884 175086
rect 268936 173120 268988 173126
rect 268936 173062 268988 173068
rect 268844 3868 268896 3874
rect 268844 3810 268896 3816
rect 268384 3324 268436 3330
rect 268384 3266 268436 3272
rect 268948 3126 268976 173062
rect 269224 172786 269252 175100
rect 269698 175086 270080 175114
rect 270158 175086 270448 175114
rect 270052 173074 270080 175086
rect 270052 173046 270356 173074
rect 269028 172780 269080 172786
rect 269028 172722 269080 172728
rect 269212 172780 269264 172786
rect 269212 172722 269264 172728
rect 270224 172780 270276 172786
rect 270224 172722 270276 172728
rect 269040 3398 269068 172722
rect 270236 4826 270264 172722
rect 270224 4820 270276 4826
rect 270224 4762 270276 4768
rect 270328 4146 270356 173046
rect 270316 4140 270368 4146
rect 270316 4082 270368 4088
rect 270420 4078 270448 175086
rect 270604 172990 270632 175100
rect 271078 175086 271552 175114
rect 271630 175086 271828 175114
rect 271524 173074 271552 175086
rect 271524 173046 271736 173074
rect 270592 172984 270644 172990
rect 270592 172926 270644 172932
rect 271604 172984 271656 172990
rect 271604 172926 271656 172932
rect 271616 7682 271644 172926
rect 271604 7676 271656 7682
rect 271604 7618 271656 7624
rect 270408 4072 270460 4078
rect 270408 4014 270460 4020
rect 271708 4010 271736 173046
rect 270500 4004 270552 4010
rect 270500 3946 270552 3952
rect 271696 4004 271748 4010
rect 271696 3946 271748 3952
rect 269028 3392 269080 3398
rect 269028 3334 269080 3340
rect 268936 3120 268988 3126
rect 268936 3062 268988 3068
rect 269304 2984 269356 2990
rect 269304 2926 269356 2932
rect 269316 480 269344 2926
rect 270512 480 270540 3946
rect 271800 3942 271828 175086
rect 272076 172990 272104 175100
rect 272550 175086 272932 175114
rect 273010 175086 273208 175114
rect 272904 173074 272932 175086
rect 272904 173046 273116 173074
rect 272064 172984 272116 172990
rect 272064 172926 272116 172932
rect 272984 172984 273036 172990
rect 272984 172926 273036 172932
rect 272996 6186 273024 172926
rect 272984 6180 273036 6186
rect 272984 6122 273036 6128
rect 271788 3936 271840 3942
rect 271788 3878 271840 3884
rect 273088 3874 273116 173046
rect 273076 3868 273128 3874
rect 273076 3810 273128 3816
rect 273180 3806 273208 175086
rect 273456 173330 273484 175100
rect 273444 173324 273496 173330
rect 273444 173266 273496 173272
rect 274376 173074 274404 175222
rect 274482 175086 274588 175114
rect 274376 173046 274496 173074
rect 274468 7614 274496 173046
rect 274456 7608 274508 7614
rect 274456 7550 274508 7556
rect 271696 3800 271748 3806
rect 271696 3742 271748 3748
rect 273168 3800 273220 3806
rect 273168 3742 273220 3748
rect 271708 480 271736 3742
rect 274560 3738 274588 175086
rect 274928 173126 274956 175100
rect 274916 173120 274968 173126
rect 274916 173062 274968 173068
rect 275388 172650 275416 175100
rect 275862 175086 275968 175114
rect 275836 173120 275888 173126
rect 275836 173062 275888 173068
rect 275376 172644 275428 172650
rect 275376 172586 275428 172592
rect 275848 8974 275876 173062
rect 275836 8968 275888 8974
rect 275836 8910 275888 8916
rect 272892 3732 272944 3738
rect 272892 3674 272944 3680
rect 274548 3732 274600 3738
rect 274548 3674 274600 3680
rect 272904 480 272932 3674
rect 275940 3670 275968 175086
rect 276400 172786 276428 175100
rect 276874 175086 277256 175114
rect 276388 172780 276440 172786
rect 276388 172722 276440 172728
rect 277124 172780 277176 172786
rect 277124 172722 277176 172728
rect 277136 15910 277164 172722
rect 277124 15904 277176 15910
rect 277124 15846 277176 15852
rect 277228 6254 277256 175086
rect 277216 6248 277268 6254
rect 277216 6190 277268 6196
rect 274088 3664 274140 3670
rect 274088 3606 274140 3612
rect 275928 3664 275980 3670
rect 275928 3606 275980 3612
rect 274100 480 274128 3606
rect 277320 3602 277348 175100
rect 277780 173126 277808 175100
rect 278254 175086 278636 175114
rect 277768 173120 277820 173126
rect 277768 173062 277820 173068
rect 278044 172644 278096 172650
rect 278044 172586 278096 172592
rect 278056 9042 278084 172586
rect 278608 13190 278636 175086
rect 278688 173120 278740 173126
rect 278688 173062 278740 173068
rect 278596 13184 278648 13190
rect 278596 13126 278648 13132
rect 278700 10402 278728 173062
rect 278792 172650 278820 175100
rect 279252 172922 279280 175100
rect 279726 175086 279924 175114
rect 279240 172916 279292 172922
rect 279240 172858 279292 172864
rect 278780 172644 278832 172650
rect 278780 172586 278832 172592
rect 279896 151094 279924 175086
rect 279976 172916 280028 172922
rect 279976 172858 280028 172864
rect 279884 151088 279936 151094
rect 279884 151030 279936 151036
rect 279988 11830 280016 172858
rect 280172 172650 280200 175100
rect 280724 173126 280752 175100
rect 281184 173262 281212 175100
rect 281172 173256 281224 173262
rect 281172 173198 281224 173204
rect 281644 173126 281672 175100
rect 280712 173120 280764 173126
rect 280712 173062 280764 173068
rect 281356 173120 281408 173126
rect 281356 173062 281408 173068
rect 281632 173120 281684 173126
rect 282472 173108 282500 175222
rect 282578 175086 282776 175114
rect 282472 173080 282684 173108
rect 281632 173062 281684 173068
rect 280068 172644 280120 172650
rect 280068 172586 280120 172592
rect 280160 172644 280212 172650
rect 280160 172586 280212 172592
rect 279976 11824 280028 11830
rect 279976 11766 280028 11772
rect 278688 10396 278740 10402
rect 278688 10338 278740 10344
rect 278044 9036 278096 9042
rect 278044 8978 278096 8984
rect 276480 3596 276532 3602
rect 276480 3538 276532 3544
rect 277308 3596 277360 3602
rect 277308 3538 277360 3544
rect 275284 3324 275336 3330
rect 275284 3266 275336 3272
rect 275296 480 275324 3266
rect 276492 480 276520 3538
rect 280080 3534 280108 172586
rect 281368 17270 281396 173062
rect 281448 172644 281500 172650
rect 281448 172586 281500 172592
rect 281356 17264 281408 17270
rect 281356 17206 281408 17212
rect 277676 3528 277728 3534
rect 277676 3470 277728 3476
rect 280068 3528 280120 3534
rect 280068 3470 280120 3476
rect 277688 480 277716 3470
rect 281460 3466 281488 172586
rect 282656 13122 282684 173080
rect 282644 13116 282696 13122
rect 282644 13058 282696 13064
rect 278872 3460 278924 3466
rect 278872 3402 278924 3408
rect 281448 3460 281500 3466
rect 281448 3402 281500 3408
rect 278884 480 278912 3402
rect 282460 3392 282512 3398
rect 282460 3334 282512 3340
rect 281264 3324 281316 3330
rect 281264 3266 281316 3272
rect 280068 3256 280120 3262
rect 280068 3198 280120 3204
rect 280080 480 280108 3198
rect 281276 480 281304 3266
rect 282472 480 282500 3334
rect 282748 2990 282776 175086
rect 282828 173120 282880 173126
rect 282828 173062 282880 173068
rect 282736 2984 282788 2990
rect 282736 2926 282788 2932
rect 282840 2854 282868 173062
rect 283116 172582 283144 175100
rect 283576 172650 283604 175100
rect 284050 175086 284156 175114
rect 283564 172644 283616 172650
rect 283564 172586 283616 172592
rect 283104 172576 283156 172582
rect 283104 172518 283156 172524
rect 283656 4820 283708 4826
rect 283656 4762 283708 4768
rect 282828 2848 282880 2854
rect 282828 2790 282880 2796
rect 283668 480 283696 4762
rect 284128 3058 284156 175086
rect 284496 172582 284524 175100
rect 284970 175086 285444 175114
rect 285522 175086 285628 175114
rect 284208 172576 284260 172582
rect 284208 172518 284260 172524
rect 284484 172576 284536 172582
rect 284484 172518 284536 172524
rect 284116 3052 284168 3058
rect 284116 2994 284168 3000
rect 284220 2922 284248 172518
rect 285416 14482 285444 175086
rect 285496 172576 285548 172582
rect 285496 172518 285548 172524
rect 285404 14476 285456 14482
rect 285404 14418 285456 14424
rect 284760 4140 284812 4146
rect 284760 4082 284812 4088
rect 284208 2916 284260 2922
rect 284208 2858 284260 2864
rect 284772 480 284800 4082
rect 285508 3126 285536 172518
rect 285600 3262 285628 175086
rect 285968 172582 285996 175100
rect 286442 175086 286824 175114
rect 285956 172576 286008 172582
rect 285956 172518 286008 172524
rect 286796 18630 286824 175086
rect 286784 18624 286836 18630
rect 286784 18566 286836 18572
rect 285956 4072 286008 4078
rect 285956 4014 286008 4020
rect 285588 3256 285640 3262
rect 285588 3198 285640 3204
rect 285496 3120 285548 3126
rect 285496 3062 285548 3068
rect 285968 480 285996 4014
rect 286888 3398 286916 175100
rect 287348 172582 287376 175100
rect 287914 175086 288296 175114
rect 287704 173324 287756 173330
rect 287704 173266 287756 173272
rect 286968 172576 287020 172582
rect 286968 172518 287020 172524
rect 287336 172576 287388 172582
rect 287336 172518 287388 172524
rect 286876 3392 286928 3398
rect 286876 3334 286928 3340
rect 286980 3194 287008 172518
rect 287152 7676 287204 7682
rect 287152 7618 287204 7624
rect 286968 3188 287020 3194
rect 286968 3130 287020 3136
rect 287164 480 287192 7618
rect 287716 5574 287744 173266
rect 288268 10334 288296 175086
rect 288360 173262 288388 175100
rect 288348 173256 288400 173262
rect 288348 173198 288400 173204
rect 288820 172582 288848 175100
rect 289294 175086 289584 175114
rect 288348 172576 288400 172582
rect 288348 172518 288400 172524
rect 288808 172576 288860 172582
rect 288808 172518 288860 172524
rect 288256 10328 288308 10334
rect 288256 10270 288308 10276
rect 287704 5568 287756 5574
rect 287704 5510 287756 5516
rect 288360 5114 288388 172518
rect 289556 11762 289584 175086
rect 289648 175086 289754 175114
rect 289544 11756 289596 11762
rect 289544 11698 289596 11704
rect 288176 5086 288388 5114
rect 288176 3330 288204 5086
rect 289648 4282 289676 175086
rect 290292 172582 290320 175100
rect 290766 175086 291056 175114
rect 290464 172644 290516 172650
rect 290464 172586 290516 172592
rect 289728 172576 289780 172582
rect 289728 172518 289780 172524
rect 290280 172576 290332 172582
rect 290280 172518 290332 172524
rect 289636 4276 289688 4282
rect 289636 4218 289688 4224
rect 289740 4146 289768 172518
rect 290476 6186 290504 172586
rect 291028 19990 291056 175086
rect 291212 172650 291240 175100
rect 291200 172644 291252 172650
rect 291200 172586 291252 172592
rect 291672 172582 291700 175100
rect 292146 175086 292344 175114
rect 291108 172576 291160 172582
rect 291108 172518 291160 172524
rect 291660 172576 291712 172582
rect 291660 172518 291712 172524
rect 291016 19984 291068 19990
rect 291016 19926 291068 19932
rect 290464 6180 290516 6186
rect 290464 6122 290516 6128
rect 290740 6044 290792 6050
rect 290740 5986 290792 5992
rect 289728 4140 289780 4146
rect 289728 4082 289780 4088
rect 288348 4004 288400 4010
rect 288348 3946 288400 3952
rect 288164 3324 288216 3330
rect 288164 3266 288216 3272
rect 288360 480 288388 3946
rect 289544 3936 289596 3942
rect 289544 3878 289596 3884
rect 289556 480 289584 3878
rect 290752 480 290780 5986
rect 291120 4078 291148 172518
rect 292316 21418 292344 175086
rect 292684 172650 292712 175100
rect 292396 172644 292448 172650
rect 292396 172586 292448 172592
rect 292672 172644 292724 172650
rect 292672 172586 292724 172592
rect 292304 21412 292356 21418
rect 292304 21354 292356 21360
rect 292408 4350 292436 172586
rect 293144 172582 293172 175100
rect 293618 175086 293724 175114
rect 292488 172576 292540 172582
rect 292488 172518 292540 172524
rect 293132 172576 293184 172582
rect 293132 172518 293184 172524
rect 292396 4344 292448 4350
rect 292396 4286 292448 4292
rect 291108 4072 291160 4078
rect 291108 4014 291160 4020
rect 292500 4010 292528 172518
rect 293696 4554 293724 175086
rect 293776 172644 293828 172650
rect 293776 172586 293828 172592
rect 293684 4548 293736 4554
rect 293684 4490 293736 4496
rect 293788 4418 293816 172586
rect 294064 172582 294092 175100
rect 294524 172650 294552 175100
rect 295090 175086 295196 175114
rect 294512 172644 294564 172650
rect 294512 172586 294564 172592
rect 293868 172576 293920 172582
rect 293868 172518 293920 172524
rect 294052 172576 294104 172582
rect 294052 172518 294104 172524
rect 295064 172576 295116 172582
rect 295064 172518 295116 172524
rect 293776 4412 293828 4418
rect 293776 4354 293828 4360
rect 292488 4004 292540 4010
rect 292488 3946 292540 3952
rect 293880 3942 293908 172518
rect 294328 5568 294380 5574
rect 294328 5510 294380 5516
rect 293868 3936 293920 3942
rect 293868 3878 293920 3884
rect 291936 3868 291988 3874
rect 291936 3810 291988 3816
rect 291948 480 291976 3810
rect 293132 3800 293184 3806
rect 293132 3742 293184 3748
rect 293144 480 293172 3742
rect 294340 480 294368 5510
rect 295076 4486 295104 172518
rect 295168 4690 295196 175086
rect 295536 172650 295564 175100
rect 295248 172644 295300 172650
rect 295248 172586 295300 172592
rect 295524 172644 295576 172650
rect 295524 172586 295576 172592
rect 295156 4684 295208 4690
rect 295156 4626 295208 4632
rect 295064 4480 295116 4486
rect 295064 4422 295116 4428
rect 295260 3874 295288 172586
rect 295996 172582 296024 175100
rect 295984 172576 296036 172582
rect 295984 172518 296036 172524
rect 295524 7608 295576 7614
rect 295524 7550 295576 7556
rect 295248 3868 295300 3874
rect 295248 3810 295300 3816
rect 295536 480 295564 7550
rect 296456 5506 296484 175100
rect 297008 172650 297036 175100
rect 296536 172644 296588 172650
rect 296536 172586 296588 172592
rect 296996 172644 297048 172650
rect 296996 172586 297048 172592
rect 296444 5500 296496 5506
rect 296444 5442 296496 5448
rect 296548 4622 296576 172586
rect 297468 172582 297496 175100
rect 297836 175086 297942 175114
rect 296628 172576 296680 172582
rect 296628 172518 296680 172524
rect 297456 172576 297508 172582
rect 297456 172518 297508 172524
rect 296536 4616 296588 4622
rect 296536 4558 296588 4564
rect 296640 3806 296668 172518
rect 297732 8968 297784 8974
rect 297732 8910 297784 8916
rect 296628 3800 296680 3806
rect 296628 3742 296680 3748
rect 296720 3732 296772 3738
rect 296720 3674 296772 3680
rect 296732 480 296760 3674
rect 297744 3482 297772 8910
rect 297836 5438 297864 175086
rect 297916 172644 297968 172650
rect 297916 172586 297968 172592
rect 297824 5432 297876 5438
rect 297824 5374 297876 5380
rect 297928 4758 297956 172586
rect 298388 172582 298416 175100
rect 298848 172650 298876 175100
rect 299308 175086 299414 175114
rect 298836 172644 298888 172650
rect 298836 172586 298888 172592
rect 298008 172576 298060 172582
rect 298008 172518 298060 172524
rect 298376 172576 298428 172582
rect 298376 172518 298428 172524
rect 299204 172576 299256 172582
rect 299204 172518 299256 172524
rect 297916 4752 297968 4758
rect 297916 4694 297968 4700
rect 298020 3738 298048 172518
rect 299112 9036 299164 9042
rect 299112 8978 299164 8984
rect 298008 3732 298060 3738
rect 298008 3674 298060 3680
rect 297744 3454 297956 3482
rect 297928 480 297956 3454
rect 299124 480 299152 8978
rect 299216 8226 299244 172518
rect 299204 8220 299256 8226
rect 299204 8162 299256 8168
rect 299308 5370 299336 175086
rect 299860 172650 299888 175100
rect 299388 172644 299440 172650
rect 299388 172586 299440 172592
rect 299848 172644 299900 172650
rect 299848 172586 299900 172592
rect 299296 5364 299348 5370
rect 299296 5306 299348 5312
rect 299400 3777 299428 172586
rect 300320 172582 300348 175100
rect 300688 175086 300794 175114
rect 300584 172644 300636 172650
rect 300584 172586 300636 172592
rect 300308 172576 300360 172582
rect 300308 172518 300360 172524
rect 300596 8158 300624 172586
rect 300584 8152 300636 8158
rect 300584 8094 300636 8100
rect 300688 5302 300716 175086
rect 301240 172582 301268 175100
rect 301806 175086 302188 175114
rect 300768 172576 300820 172582
rect 300768 172518 300820 172524
rect 301228 172576 301280 172582
rect 301228 172518 301280 172524
rect 302056 172576 302108 172582
rect 302056 172518 302108 172524
rect 300676 5296 300728 5302
rect 300676 5238 300728 5244
rect 299386 3768 299442 3777
rect 300780 3738 300808 172518
rect 300860 15904 300912 15910
rect 300860 15846 300912 15852
rect 299386 3703 299442 3712
rect 300768 3732 300820 3738
rect 300768 3674 300820 3680
rect 300308 3664 300360 3670
rect 300308 3606 300360 3612
rect 300320 480 300348 3606
rect 300872 610 300900 15846
rect 302068 8090 302096 172518
rect 302056 8084 302108 8090
rect 302056 8026 302108 8032
rect 302160 3641 302188 175086
rect 302252 172582 302280 175100
rect 302712 172650 302740 175100
rect 303186 175086 303568 175114
rect 302700 172644 302752 172650
rect 302700 172586 302752 172592
rect 303344 172644 303396 172650
rect 303344 172586 303396 172592
rect 302240 172576 302292 172582
rect 302240 172518 302292 172524
rect 303356 8022 303384 172586
rect 303436 172576 303488 172582
rect 303436 172518 303488 172524
rect 303344 8016 303396 8022
rect 303344 7958 303396 7964
rect 302608 6248 302660 6254
rect 302608 6190 302660 6196
rect 302146 3632 302202 3641
rect 302146 3567 302202 3576
rect 300860 604 300912 610
rect 300860 546 300912 552
rect 301412 604 301464 610
rect 301412 546 301464 552
rect 301424 480 301452 546
rect 302620 480 302648 6190
rect 303448 5234 303476 172518
rect 303436 5228 303488 5234
rect 303436 5170 303488 5176
rect 303540 3505 303568 175086
rect 303632 172582 303660 175100
rect 303620 172576 303672 172582
rect 303620 172518 303672 172524
rect 304552 171034 304580 175222
rect 304658 175086 304948 175114
rect 304816 172576 304868 172582
rect 304816 172518 304868 172524
rect 304552 171006 304764 171034
rect 304736 7954 304764 171006
rect 304724 7948 304776 7954
rect 304724 7890 304776 7896
rect 304828 5166 304856 172518
rect 304816 5160 304868 5166
rect 304816 5102 304868 5108
rect 304920 3602 304948 175086
rect 305104 172582 305132 175100
rect 305564 172650 305592 175100
rect 306038 175086 306328 175114
rect 305552 172644 305604 172650
rect 305552 172586 305604 172592
rect 306104 172644 306156 172650
rect 306104 172586 306156 172592
rect 305092 172576 305144 172582
rect 305092 172518 305144 172524
rect 305000 13184 305052 13190
rect 305000 13126 305052 13132
rect 305012 3738 305040 13126
rect 305092 10396 305144 10402
rect 305092 10338 305144 10344
rect 305000 3732 305052 3738
rect 305000 3674 305052 3680
rect 303804 3596 303856 3602
rect 303804 3538 303856 3544
rect 304908 3596 304960 3602
rect 304908 3538 304960 3544
rect 303526 3496 303582 3505
rect 303526 3431 303582 3440
rect 303816 480 303844 3538
rect 305104 3482 305132 10338
rect 306116 7886 306144 172586
rect 306196 172576 306248 172582
rect 306196 172518 306248 172524
rect 306104 7880 306156 7886
rect 306104 7822 306156 7828
rect 306208 5098 306236 172518
rect 306196 5092 306248 5098
rect 306196 5034 306248 5040
rect 306104 3732 306156 3738
rect 306104 3674 306156 3680
rect 305012 3454 305132 3482
rect 306116 3482 306144 3674
rect 306116 3454 306236 3482
rect 305012 480 305040 3454
rect 306208 480 306236 3454
rect 306300 3369 306328 175086
rect 306576 172582 306604 175100
rect 307036 172650 307064 175100
rect 307496 172922 307524 175100
rect 307484 172916 307536 172922
rect 307484 172858 307536 172864
rect 307024 172644 307076 172650
rect 307024 172586 307076 172592
rect 307576 172644 307628 172650
rect 307576 172586 307628 172592
rect 306564 172576 306616 172582
rect 306564 172518 306616 172524
rect 307588 7818 307616 172586
rect 307956 172582 307984 175100
rect 308430 175086 308904 175114
rect 308982 175086 309088 175114
rect 307668 172576 307720 172582
rect 307668 172518 307720 172524
rect 307944 172576 307996 172582
rect 307944 172518 307996 172524
rect 307576 7812 307628 7818
rect 307576 7754 307628 7760
rect 307680 5030 307708 172518
rect 307760 11824 307812 11830
rect 307760 11766 307812 11772
rect 307668 5024 307720 5030
rect 307668 4966 307720 4972
rect 307392 3528 307444 3534
rect 307392 3470 307444 3476
rect 306286 3360 306342 3369
rect 306286 3295 306342 3304
rect 307404 480 307432 3470
rect 307772 610 307800 11766
rect 308876 7750 308904 175086
rect 308956 172576 309008 172582
rect 308956 172518 309008 172524
rect 308864 7744 308916 7750
rect 308864 7686 308916 7692
rect 308968 4962 308996 172518
rect 308956 4956 309008 4962
rect 308956 4898 309008 4904
rect 309060 3534 309088 175086
rect 309428 172582 309456 175100
rect 309416 172576 309468 172582
rect 309416 172518 309468 172524
rect 310256 171034 310284 175222
rect 310348 172990 310376 175100
rect 310336 172984 310388 172990
rect 310336 172926 310388 172932
rect 310808 172582 310836 175100
rect 311374 175086 311664 175114
rect 310428 172576 310480 172582
rect 310428 172518 310480 172524
rect 310796 172576 310848 172582
rect 310796 172518 310848 172524
rect 310256 171006 310376 171034
rect 309140 151088 309192 151094
rect 309140 151030 309192 151036
rect 309048 3528 309100 3534
rect 309048 3470 309100 3476
rect 309152 610 309180 151030
rect 310348 7682 310376 171006
rect 310336 7676 310388 7682
rect 310336 7618 310388 7624
rect 310440 4894 310468 172518
rect 311636 7614 311664 175086
rect 311716 172576 311768 172582
rect 311716 172518 311768 172524
rect 311624 7608 311676 7614
rect 311624 7550 311676 7556
rect 310428 4888 310480 4894
rect 310428 4830 310480 4836
rect 311728 4826 311756 172518
rect 311716 4820 311768 4826
rect 311716 4762 311768 4768
rect 311820 3466 311848 175100
rect 312280 170406 312308 175100
rect 312754 175086 313228 175114
rect 312544 173392 312596 173398
rect 312544 173334 312596 173340
rect 312268 170400 312320 170406
rect 312268 170342 312320 170348
rect 311900 17264 311952 17270
rect 311900 17206 311952 17212
rect 310980 3460 311032 3466
rect 310980 3402 311032 3408
rect 311808 3460 311860 3466
rect 311808 3402 311860 3408
rect 307760 604 307812 610
rect 307760 546 307812 552
rect 308588 604 308640 610
rect 308588 546 308640 552
rect 309140 604 309192 610
rect 309140 546 309192 552
rect 309784 604 309836 610
rect 309784 546 309836 552
rect 308600 480 308628 546
rect 309796 480 309824 546
rect 310992 480 311020 3402
rect 311912 626 311940 17206
rect 312556 9654 312584 173334
rect 312544 9648 312596 9654
rect 312544 9590 312596 9596
rect 313200 7070 313228 175086
rect 313292 172582 313320 175100
rect 313766 175086 314056 175114
rect 314226 175086 314516 175114
rect 313280 172576 313332 172582
rect 313280 172518 313332 172524
rect 314028 171034 314056 175086
rect 314028 171006 314424 171034
rect 314396 156738 314424 171006
rect 314384 156732 314436 156738
rect 314384 156674 314436 156680
rect 313372 9648 313424 9654
rect 313372 9590 313424 9596
rect 313188 7064 313240 7070
rect 313188 7006 313240 7012
rect 311912 598 312216 626
rect 312188 480 312216 598
rect 313384 480 313412 9590
rect 314488 7138 314516 175086
rect 314672 173058 314700 175100
rect 314660 173052 314712 173058
rect 314660 172994 314712 173000
rect 315132 172582 315160 175100
rect 315698 175086 315988 175114
rect 314568 172576 314620 172582
rect 314568 172518 314620 172524
rect 315120 172576 315172 172582
rect 315120 172518 315172 172524
rect 315856 172576 315908 172582
rect 315856 172518 315908 172524
rect 314476 7132 314528 7138
rect 314476 7074 314528 7080
rect 314580 2938 314608 172518
rect 315868 155310 315896 172518
rect 315856 155304 315908 155310
rect 315856 155246 315908 155252
rect 314660 13116 314712 13122
rect 314660 13058 314712 13064
rect 314672 3074 314700 13058
rect 315960 8498 315988 175086
rect 316144 172582 316172 175100
rect 316618 175086 316908 175114
rect 317078 175086 317276 175114
rect 316132 172576 316184 172582
rect 316132 172518 316184 172524
rect 316880 171034 316908 175086
rect 316880 171006 317184 171034
rect 317156 153950 317184 171006
rect 317144 153944 317196 153950
rect 317144 153886 317196 153892
rect 317248 8566 317276 175086
rect 317524 173262 317552 175100
rect 318090 175086 318380 175114
rect 318550 175086 318748 175114
rect 317512 173256 317564 173262
rect 317512 173198 317564 173204
rect 317328 172576 317380 172582
rect 317328 172518 317380 172524
rect 317236 8560 317288 8566
rect 317236 8502 317288 8508
rect 315948 8492 316000 8498
rect 315948 8434 316000 8440
rect 314672 3046 314792 3074
rect 314580 2910 314700 2938
rect 314672 2854 314700 2910
rect 314568 2848 314620 2854
rect 314568 2790 314620 2796
rect 314660 2848 314712 2854
rect 314660 2790 314712 2796
rect 314580 480 314608 2790
rect 314764 610 314792 3046
rect 317340 2990 317368 172518
rect 318352 171034 318380 175086
rect 318352 171006 318656 171034
rect 318628 152590 318656 171006
rect 318616 152584 318668 152590
rect 318616 152526 318668 152532
rect 318720 8634 318748 175086
rect 318996 172582 319024 175100
rect 318984 172576 319036 172582
rect 318984 172518 319036 172524
rect 319824 171034 319852 175222
rect 319930 175086 320036 175114
rect 319824 171006 319944 171034
rect 319916 151162 319944 171006
rect 319904 151156 319956 151162
rect 319904 151098 319956 151104
rect 320008 8702 320036 175086
rect 320468 173874 320496 175100
rect 320456 173868 320508 173874
rect 320456 173810 320508 173816
rect 320088 172576 320140 172582
rect 320088 172518 320140 172524
rect 319996 8696 320048 8702
rect 319996 8638 320048 8644
rect 318708 8628 318760 8634
rect 318708 8570 318760 8576
rect 319260 6180 319312 6186
rect 319260 6122 319312 6128
rect 316960 2984 317012 2990
rect 316960 2926 317012 2932
rect 317328 2984 317380 2990
rect 317328 2926 317380 2932
rect 314752 604 314804 610
rect 314752 546 314804 552
rect 315764 604 315816 610
rect 315764 546 315816 552
rect 315776 480 315804 546
rect 316972 480 317000 2926
rect 318064 2916 318116 2922
rect 318064 2858 318116 2864
rect 318076 480 318104 2858
rect 319272 480 319300 6122
rect 320100 2922 320128 172518
rect 321296 171034 321324 175222
rect 321402 175086 321508 175114
rect 321296 171006 321416 171034
rect 321388 149802 321416 171006
rect 321376 149796 321428 149802
rect 321376 149738 321428 149744
rect 321480 8770 321508 175086
rect 321848 172786 321876 175100
rect 322322 175086 322704 175114
rect 321836 172780 321888 172786
rect 321836 172722 321888 172728
rect 322676 148442 322704 175086
rect 322768 175086 322874 175114
rect 322664 148436 322716 148442
rect 322664 148378 322716 148384
rect 321652 14476 321704 14482
rect 321652 14418 321704 14424
rect 321468 8764 321520 8770
rect 321468 8706 321520 8712
rect 321664 3262 321692 14418
rect 322768 8838 322796 175086
rect 323320 173806 323348 175100
rect 323794 175086 324176 175114
rect 323308 173800 323360 173806
rect 323308 173742 323360 173748
rect 322848 172780 322900 172786
rect 322848 172722 322900 172728
rect 322756 8832 322808 8838
rect 322756 8774 322808 8780
rect 322860 4978 322888 172722
rect 324148 147014 324176 175086
rect 324136 147008 324188 147014
rect 324136 146950 324188 146956
rect 324240 8906 324268 175100
rect 324700 173262 324728 175100
rect 325266 175086 325556 175114
rect 324688 173256 324740 173262
rect 324688 173198 324740 173204
rect 324228 8900 324280 8906
rect 324228 8842 324280 8848
rect 325528 5642 325556 175086
rect 325712 173262 325740 175100
rect 326172 173738 326200 175100
rect 326646 175086 327028 175114
rect 326160 173732 326212 173738
rect 326160 173674 326212 173680
rect 325608 173256 325660 173262
rect 325608 173198 325660 173204
rect 325700 173256 325752 173262
rect 325700 173198 325752 173204
rect 326896 173256 326948 173262
rect 326896 173198 326948 173204
rect 325516 5636 325568 5642
rect 325516 5578 325568 5584
rect 322768 4950 322888 4978
rect 321652 3256 321704 3262
rect 321652 3198 321704 3204
rect 321652 3120 321704 3126
rect 321652 3062 321704 3068
rect 320456 3052 320508 3058
rect 320456 2994 320508 3000
rect 320088 2916 320140 2922
rect 320088 2858 320140 2864
rect 320468 480 320496 2994
rect 321664 480 321692 3062
rect 322768 3058 322796 4950
rect 322848 3256 322900 3262
rect 322848 3198 322900 3204
rect 322756 3052 322808 3058
rect 322756 2994 322808 3000
rect 322860 480 322888 3198
rect 324044 3188 324096 3194
rect 324044 3130 324096 3136
rect 324056 480 324084 3130
rect 325620 3126 325648 173198
rect 325700 18624 325752 18630
rect 325700 18566 325752 18572
rect 325608 3120 325660 3126
rect 325608 3062 325660 3068
rect 325240 2984 325292 2990
rect 325240 2926 325292 2932
rect 325252 480 325280 2926
rect 325712 610 325740 18566
rect 326908 9654 326936 173198
rect 326896 9648 326948 9654
rect 326896 9590 326948 9596
rect 327000 5710 327028 175086
rect 327092 172650 327120 175100
rect 327644 173194 327672 175100
rect 328118 175086 328316 175114
rect 327632 173188 327684 173194
rect 327632 173130 327684 173136
rect 327080 172644 327132 172650
rect 327080 172586 327132 172592
rect 328184 172644 328236 172650
rect 328184 172586 328236 172592
rect 328196 9586 328224 172586
rect 328184 9580 328236 9586
rect 328184 9522 328236 9528
rect 328288 5778 328316 175086
rect 328564 173194 328592 175100
rect 329024 173670 329052 175100
rect 329590 175086 329788 175114
rect 329012 173664 329064 173670
rect 329012 173606 329064 173612
rect 328368 173188 328420 173194
rect 328368 173130 328420 173136
rect 328552 173188 328604 173194
rect 328552 173130 328604 173136
rect 329656 173188 329708 173194
rect 329656 173130 329708 173136
rect 328276 5772 328328 5778
rect 328276 5714 328328 5720
rect 326988 5704 327040 5710
rect 326988 5646 327040 5652
rect 327632 3392 327684 3398
rect 327632 3334 327684 3340
rect 325700 604 325752 610
rect 325700 546 325752 552
rect 326436 604 326488 610
rect 326436 546 326488 552
rect 326448 480 326476 546
rect 327644 480 327672 3334
rect 328380 3194 328408 173130
rect 329668 9518 329696 173130
rect 329656 9512 329708 9518
rect 329656 9454 329708 9460
rect 329760 5846 329788 175086
rect 330036 173194 330064 175100
rect 330496 173262 330524 175100
rect 330970 175086 331076 175114
rect 330484 173256 330536 173262
rect 330484 173198 330536 173204
rect 330024 173188 330076 173194
rect 330024 173130 330076 173136
rect 330944 173188 330996 173194
rect 330944 173130 330996 173136
rect 329840 10328 329892 10334
rect 329840 10270 329892 10276
rect 329748 5840 329800 5846
rect 329748 5782 329800 5788
rect 328828 3324 328880 3330
rect 328828 3266 328880 3272
rect 328368 3188 328420 3194
rect 328368 3130 328420 3136
rect 328840 480 328868 3266
rect 329852 626 329880 10270
rect 330956 9450 330984 173130
rect 330944 9444 330996 9450
rect 330944 9386 330996 9392
rect 331048 5914 331076 175086
rect 331312 173324 331364 173330
rect 331312 173266 331364 173272
rect 331128 173256 331180 173262
rect 331128 173198 331180 173204
rect 331036 5908 331088 5914
rect 331036 5850 331088 5856
rect 331140 3262 331168 173198
rect 331128 3256 331180 3262
rect 331128 3198 331180 3204
rect 331324 626 331352 173266
rect 331416 173194 331444 175100
rect 331968 173602 331996 175100
rect 332442 175086 332548 175114
rect 331956 173596 332008 173602
rect 331956 173538 332008 173544
rect 331404 173188 331456 173194
rect 331404 173130 331456 173136
rect 332416 173188 332468 173194
rect 332416 173130 332468 173136
rect 332428 9382 332456 173130
rect 332416 9376 332468 9382
rect 332416 9318 332468 9324
rect 332520 5982 332548 175086
rect 332888 173194 332916 175100
rect 333348 173262 333376 175100
rect 333336 173256 333388 173262
rect 333336 173198 333388 173204
rect 332876 173188 332928 173194
rect 332876 173130 332928 173136
rect 333704 173188 333756 173194
rect 333704 173130 333756 173136
rect 332600 11756 332652 11762
rect 332600 11698 332652 11704
rect 332508 5976 332560 5982
rect 332508 5918 332560 5924
rect 332416 4140 332468 4146
rect 332416 4082 332468 4088
rect 329852 598 330064 626
rect 330036 480 330064 598
rect 331232 598 331352 626
rect 331232 480 331260 598
rect 332428 480 332456 4082
rect 332612 610 332640 11698
rect 333716 9314 333744 173130
rect 333704 9308 333756 9314
rect 333704 9250 333756 9256
rect 333808 6050 333836 175100
rect 333888 173256 333940 173262
rect 333888 173198 333940 173204
rect 333796 6044 333848 6050
rect 333796 5986 333848 5992
rect 333900 3330 333928 173198
rect 334360 172650 334388 175100
rect 334820 173534 334848 175100
rect 334808 173528 334860 173534
rect 334808 173470 334860 173476
rect 334348 172644 334400 172650
rect 334348 172586 334400 172592
rect 335176 172644 335228 172650
rect 335176 172586 335228 172592
rect 335188 9246 335216 172586
rect 335176 9240 335228 9246
rect 335176 9182 335228 9188
rect 335280 6118 335308 175100
rect 335740 173194 335768 175100
rect 336214 175086 336688 175114
rect 335728 173188 335780 173194
rect 335728 173130 335780 173136
rect 336556 173188 336608 173194
rect 336556 173130 336608 173136
rect 336568 9178 336596 173130
rect 336556 9172 336608 9178
rect 336556 9114 336608 9120
rect 335268 6112 335320 6118
rect 335268 6054 335320 6060
rect 334716 4276 334768 4282
rect 334716 4218 334768 4224
rect 333888 3324 333940 3330
rect 333888 3266 333940 3272
rect 332600 604 332652 610
rect 332600 546 332652 552
rect 333612 604 333664 610
rect 333612 546 333664 552
rect 333624 480 333652 546
rect 334728 480 334756 4218
rect 335912 4072 335964 4078
rect 335912 4014 335964 4020
rect 335924 480 335952 4014
rect 336660 3398 336688 175086
rect 336752 173194 336780 175100
rect 337212 173262 337240 175100
rect 337672 173466 337700 175100
rect 337660 173460 337712 173466
rect 337660 173402 337712 173408
rect 337200 173256 337252 173262
rect 337200 173198 337252 173204
rect 337936 173256 337988 173262
rect 337936 173198 337988 173204
rect 336740 173188 336792 173194
rect 336740 173130 336792 173136
rect 336740 19984 336792 19990
rect 336740 19926 336792 19932
rect 336648 3392 336700 3398
rect 336648 3334 336700 3340
rect 336752 610 336780 19926
rect 337948 9110 337976 173198
rect 338132 173194 338160 175100
rect 338592 173262 338620 175100
rect 339158 175086 339448 175114
rect 338580 173256 338632 173262
rect 338580 173198 338632 173204
rect 339224 173256 339276 173262
rect 339224 173198 339276 173204
rect 338028 173188 338080 173194
rect 338028 173130 338080 173136
rect 338120 173188 338172 173194
rect 338120 173130 338172 173136
rect 337936 9104 337988 9110
rect 337936 9046 337988 9052
rect 338040 6866 338068 173130
rect 339236 9042 339264 173198
rect 339316 173188 339368 173194
rect 339316 173130 339368 173136
rect 339224 9036 339276 9042
rect 339224 8978 339276 8984
rect 338028 6860 338080 6866
rect 338028 6802 338080 6808
rect 339328 6798 339356 173130
rect 339316 6792 339368 6798
rect 339316 6734 339368 6740
rect 338304 4344 338356 4350
rect 338304 4286 338356 4292
rect 336740 604 336792 610
rect 336740 546 336792 552
rect 337108 604 337160 610
rect 337108 546 337160 552
rect 337120 480 337148 546
rect 338316 480 338344 4286
rect 339420 4146 339448 175086
rect 339604 173194 339632 175100
rect 340064 173262 340092 175100
rect 340524 173398 340552 175100
rect 340512 173392 340564 173398
rect 340512 173334 340564 173340
rect 340052 173256 340104 173262
rect 340052 173198 340104 173204
rect 340696 173256 340748 173262
rect 340696 173198 340748 173204
rect 339592 173188 339644 173194
rect 339592 173130 339644 173136
rect 339592 21412 339644 21418
rect 339592 21354 339644 21360
rect 339408 4140 339460 4146
rect 339408 4082 339460 4088
rect 339500 4004 339552 4010
rect 339500 3946 339552 3952
rect 339512 480 339540 3946
rect 339604 610 339632 21354
rect 340708 8974 340736 173198
rect 340788 173188 340840 173194
rect 340788 173130 340840 173136
rect 340696 8968 340748 8974
rect 340696 8910 340748 8916
rect 340800 6730 340828 173130
rect 340984 172786 341012 175100
rect 341904 173074 341932 175222
rect 342010 175086 342208 175114
rect 341904 173046 342024 173074
rect 340972 172780 341024 172786
rect 340972 172722 341024 172728
rect 341996 137290 342024 173046
rect 342076 172780 342128 172786
rect 342076 172722 342128 172728
rect 341984 137284 342036 137290
rect 341984 137226 342036 137232
rect 340788 6724 340840 6730
rect 340788 6666 340840 6672
rect 342088 6662 342116 172722
rect 342076 6656 342128 6662
rect 342076 6598 342128 6604
rect 341892 4412 341944 4418
rect 341892 4354 341944 4360
rect 339592 604 339644 610
rect 339592 546 339644 552
rect 340696 604 340748 610
rect 340696 546 340748 552
rect 340708 480 340736 546
rect 341904 480 341932 4354
rect 342180 4078 342208 175086
rect 342456 173194 342484 175100
rect 342444 173188 342496 173194
rect 342444 173130 342496 173136
rect 343376 173074 343404 175222
rect 352116 175222 352498 175250
rect 353588 175222 353970 175250
rect 362158 175222 362540 175250
rect 377430 175222 377812 175250
rect 343468 173330 343496 175100
rect 343456 173324 343508 173330
rect 343456 173266 343508 173272
rect 343928 173194 343956 175100
rect 344402 175086 344784 175114
rect 344862 175086 344968 175114
rect 343548 173188 343600 173194
rect 343548 173130 343600 173136
rect 343916 173188 343968 173194
rect 343916 173130 343968 173136
rect 343376 173046 343496 173074
rect 343468 133210 343496 173046
rect 343456 133204 343508 133210
rect 343456 133146 343508 133152
rect 343560 6594 343588 173130
rect 344756 135930 344784 175086
rect 344836 173188 344888 173194
rect 344836 173130 344888 173136
rect 344744 135924 344796 135930
rect 344744 135866 344796 135872
rect 343548 6588 343600 6594
rect 343548 6530 343600 6536
rect 344848 6526 344876 173130
rect 344836 6520 344888 6526
rect 344836 6462 344888 6468
rect 344284 4548 344336 4554
rect 344284 4490 344336 4496
rect 342168 4072 342220 4078
rect 342168 4014 342220 4020
rect 343088 3936 343140 3942
rect 343088 3878 343140 3884
rect 343100 480 343128 3878
rect 344296 480 344324 4490
rect 344940 4010 344968 175086
rect 345308 173194 345336 175100
rect 345874 175086 346256 175114
rect 345296 173188 345348 173194
rect 345296 173130 345348 173136
rect 346228 130422 346256 175086
rect 346320 173346 346348 175100
rect 346320 173318 346440 173346
rect 346308 173188 346360 173194
rect 346308 173130 346360 173136
rect 346216 130416 346268 130422
rect 346216 130358 346268 130364
rect 346320 6458 346348 173130
rect 346412 172854 346440 173318
rect 346780 173194 346808 175100
rect 347254 175086 347544 175114
rect 346768 173188 346820 173194
rect 346768 173130 346820 173136
rect 346400 172848 346452 172854
rect 346400 172790 346452 172796
rect 347516 131782 347544 175086
rect 347596 173188 347648 173194
rect 347596 173130 347648 173136
rect 347504 131776 347556 131782
rect 347504 131718 347556 131724
rect 346308 6452 346360 6458
rect 346308 6394 346360 6400
rect 347608 6390 347636 173130
rect 347596 6384 347648 6390
rect 347596 6326 347648 6332
rect 345480 4480 345532 4486
rect 345480 4422 345532 4428
rect 344928 4004 344980 4010
rect 344928 3946 344980 3952
rect 345492 480 345520 4422
rect 347700 3942 347728 175100
rect 348252 173194 348280 175100
rect 348726 175086 349016 175114
rect 348240 173188 348292 173194
rect 348240 173130 348292 173136
rect 348988 127634 349016 175086
rect 349172 173262 349200 175100
rect 349160 173256 349212 173262
rect 349160 173198 349212 173204
rect 349068 173188 349120 173194
rect 349068 173130 349120 173136
rect 348976 127628 349028 127634
rect 348976 127570 349028 127576
rect 349080 6322 349108 173130
rect 349632 171834 349660 175100
rect 350106 175086 350396 175114
rect 349620 171828 349672 171834
rect 349620 171770 349672 171776
rect 349068 6316 349120 6322
rect 349068 6258 349120 6264
rect 350368 6254 350396 175086
rect 350644 173194 350672 175100
rect 350828 175086 351118 175114
rect 351578 175086 351868 175114
rect 350632 173188 350684 173194
rect 350632 173130 350684 173136
rect 350828 173074 350856 175086
rect 351736 173188 351788 173194
rect 351736 173130 351788 173136
rect 350644 173046 350856 173074
rect 350644 169046 350672 173046
rect 350632 169040 350684 169046
rect 350632 168982 350684 168988
rect 351748 11762 351776 173130
rect 351736 11756 351788 11762
rect 351736 11698 351788 11704
rect 350356 6248 350408 6254
rect 350356 6190 350408 6196
rect 351840 6186 351868 175086
rect 352024 173194 352052 175100
rect 352012 173188 352064 173194
rect 352012 173130 352064 173136
rect 352116 173074 352144 175222
rect 353050 175086 353156 175114
rect 352024 173046 352144 173074
rect 352024 167686 352052 173046
rect 352012 167680 352064 167686
rect 352012 167622 352064 167628
rect 353128 145586 353156 175086
rect 353208 173188 353260 173194
rect 353208 173130 353260 173136
rect 353116 145580 353168 145586
rect 353116 145522 353168 145528
rect 353220 10334 353248 173130
rect 353496 172786 353524 175100
rect 353484 172780 353536 172786
rect 353484 172722 353536 172728
rect 353588 172666 353616 175222
rect 354430 175086 354628 175114
rect 354496 172780 354548 172786
rect 354496 172722 354548 172728
rect 353404 172638 353616 172666
rect 353404 166326 353432 172638
rect 353392 166320 353444 166326
rect 353392 166262 353444 166268
rect 354508 129062 354536 172722
rect 354496 129056 354548 129062
rect 354496 128998 354548 129004
rect 354600 14482 354628 175086
rect 354876 172854 354904 175100
rect 354864 172848 354916 172854
rect 354864 172790 354916 172796
rect 355428 172786 355456 175100
rect 354772 172780 354824 172786
rect 354772 172722 354824 172728
rect 355416 172780 355468 172786
rect 355416 172722 355468 172728
rect 354784 164898 354812 172722
rect 354772 164892 354824 164898
rect 354772 164834 354824 164840
rect 355888 141438 355916 175100
rect 356348 172854 356376 175100
rect 356822 175086 357204 175114
rect 355968 172848 356020 172854
rect 355968 172790 356020 172796
rect 356336 172848 356388 172854
rect 356336 172790 356388 172796
rect 355876 141432 355928 141438
rect 355876 141374 355928 141380
rect 354588 14476 354640 14482
rect 354588 14418 354640 14424
rect 355980 13122 356008 172790
rect 357176 163538 357204 175086
rect 357164 163532 357216 163538
rect 357164 163474 357216 163480
rect 357268 142866 357296 175100
rect 357820 172854 357848 175100
rect 358294 175086 358584 175114
rect 357348 172848 357400 172854
rect 357348 172790 357400 172796
rect 357808 172848 357860 172854
rect 357808 172790 357860 172796
rect 357256 142860 357308 142866
rect 357256 142802 357308 142808
rect 357360 15910 357388 172790
rect 358556 162178 358584 175086
rect 358648 175086 358754 175114
rect 358544 162172 358596 162178
rect 358544 162114 358596 162120
rect 358648 144226 358676 175086
rect 359200 172854 359228 175100
rect 359766 175086 360056 175114
rect 358728 172848 358780 172854
rect 358728 172790 358780 172796
rect 359188 172848 359240 172854
rect 359188 172790 359240 172796
rect 358636 144220 358688 144226
rect 358636 144162 358688 144168
rect 358740 17270 358768 172790
rect 360028 160750 360056 175086
rect 360108 172848 360160 172854
rect 360108 172790 360160 172796
rect 360016 160744 360068 160750
rect 360016 160686 360068 160692
rect 360120 18630 360148 172790
rect 360212 172786 360240 175100
rect 360672 172854 360700 175100
rect 361146 175086 361344 175114
rect 360660 172848 360712 172854
rect 360660 172790 360712 172796
rect 360200 172780 360252 172786
rect 360200 172722 360252 172728
rect 361316 159390 361344 175086
rect 361592 172854 361620 175100
rect 362512 173074 362540 175222
rect 362618 175086 362908 175114
rect 362512 173046 362724 173074
rect 361488 172848 361540 172854
rect 361488 172790 361540 172796
rect 361580 172848 361632 172854
rect 361580 172790 361632 172796
rect 361396 172780 361448 172786
rect 361396 172722 361448 172728
rect 361304 159384 361356 159390
rect 361304 159326 361356 159332
rect 361408 138718 361436 172722
rect 361396 138712 361448 138718
rect 361396 138654 361448 138660
rect 361500 19990 361528 172790
rect 362696 153882 362724 173046
rect 362776 172848 362828 172854
rect 362776 172790 362828 172796
rect 362684 153876 362736 153882
rect 362684 153818 362736 153824
rect 362788 140078 362816 172790
rect 362776 140072 362828 140078
rect 362776 140014 362828 140020
rect 361488 19984 361540 19990
rect 361488 19926 361540 19932
rect 360108 18624 360160 18630
rect 360108 18566 360160 18572
rect 358728 17264 358780 17270
rect 358728 17206 358780 17212
rect 357348 15904 357400 15910
rect 357348 15846 357400 15852
rect 355968 13116 356020 13122
rect 355968 13058 356020 13064
rect 353208 10328 353260 10334
rect 353208 10270 353260 10276
rect 356152 8220 356204 8226
rect 356152 8162 356204 8168
rect 351828 6180 351880 6186
rect 351828 6122 351880 6128
rect 351368 5500 351420 5506
rect 351368 5442 351420 5448
rect 347872 4684 347924 4690
rect 347872 4626 347924 4632
rect 347688 3936 347740 3942
rect 347688 3878 347740 3884
rect 346676 3868 346728 3874
rect 346676 3810 346728 3816
rect 346688 480 346716 3810
rect 347884 480 347912 4626
rect 349068 4616 349120 4622
rect 349068 4558 349120 4564
rect 349080 480 349108 4558
rect 350264 3800 350316 3806
rect 350264 3742 350316 3748
rect 350276 480 350304 3742
rect 351380 480 351408 5442
rect 354956 5432 355008 5438
rect 354956 5374 355008 5380
rect 352564 4752 352616 4758
rect 352564 4694 352616 4700
rect 352576 480 352604 4694
rect 353760 3732 353812 3738
rect 353760 3674 353812 3680
rect 353772 480 353800 3674
rect 354968 480 354996 5374
rect 356164 480 356192 8162
rect 359740 8152 359792 8158
rect 359740 8094 359792 8100
rect 358544 5364 358596 5370
rect 358544 5306 358596 5312
rect 357346 3768 357402 3777
rect 357346 3703 357402 3712
rect 357360 480 357388 3703
rect 358556 480 358584 5306
rect 359752 480 359780 8094
rect 362132 5296 362184 5302
rect 362132 5238 362184 5244
rect 360936 3664 360988 3670
rect 360936 3606 360988 3612
rect 360948 480 360976 3606
rect 362144 480 362172 5238
rect 362880 4282 362908 175086
rect 363064 172854 363092 175100
rect 363538 175086 363920 175114
rect 363998 175086 364288 175114
rect 363892 173074 363920 175086
rect 363892 173046 364196 173074
rect 363052 172848 363104 172854
rect 363052 172790 363104 172796
rect 364064 172848 364116 172854
rect 364064 172790 364116 172796
rect 364076 156670 364104 172790
rect 364064 156664 364116 156670
rect 364064 156606 364116 156612
rect 364168 124914 364196 173046
rect 364156 124908 364208 124914
rect 364156 124850 364208 124856
rect 363328 8084 363380 8090
rect 363328 8026 363380 8032
rect 362868 4276 362920 4282
rect 362868 4218 362920 4224
rect 363340 480 363368 8026
rect 364260 4350 364288 175086
rect 364536 172854 364564 175100
rect 365010 175086 365392 175114
rect 365470 175086 365668 175114
rect 365364 173074 365392 175086
rect 365364 173046 365576 173074
rect 364524 172848 364576 172854
rect 364524 172790 364576 172796
rect 365444 172848 365496 172854
rect 365444 172790 365496 172796
rect 365456 155242 365484 172790
rect 365444 155236 365496 155242
rect 365444 155178 365496 155184
rect 365548 21418 365576 173046
rect 365536 21412 365588 21418
rect 365536 21354 365588 21360
rect 365640 4418 365668 175086
rect 365916 172854 365944 175100
rect 366390 175086 366864 175114
rect 366942 175086 367048 175114
rect 365904 172848 365956 172854
rect 365904 172790 365956 172796
rect 366836 152522 366864 175086
rect 366916 172848 366968 172854
rect 366916 172790 366968 172796
rect 366824 152516 366876 152522
rect 366824 152458 366876 152464
rect 366928 11914 366956 172790
rect 366836 11886 366956 11914
rect 366836 7206 366864 11886
rect 366916 8016 366968 8022
rect 366916 7958 366968 7964
rect 366824 7200 366876 7206
rect 366824 7142 366876 7148
rect 365720 5228 365772 5234
rect 365720 5170 365772 5176
rect 365628 4412 365680 4418
rect 365628 4354 365680 4360
rect 364248 4344 364300 4350
rect 364248 4286 364300 4292
rect 364522 3632 364578 3641
rect 364522 3567 364578 3576
rect 364536 480 364564 3567
rect 365732 480 365760 5170
rect 366928 480 366956 7958
rect 367020 4486 367048 175086
rect 367388 172854 367416 175100
rect 367862 175086 368244 175114
rect 368322 175086 368428 175114
rect 367376 172848 367428 172854
rect 367376 172790 367428 172796
rect 368216 151094 368244 175086
rect 368296 172848 368348 172854
rect 368296 172790 368348 172796
rect 368204 151088 368256 151094
rect 368204 151030 368256 151036
rect 368308 7274 368336 172790
rect 368296 7268 368348 7274
rect 368296 7210 368348 7216
rect 368400 4554 368428 175086
rect 368768 172854 368796 175100
rect 369334 175086 369624 175114
rect 368756 172848 368808 172854
rect 368756 172790 368808 172796
rect 369596 149734 369624 175086
rect 369676 172848 369728 172854
rect 369676 172790 369728 172796
rect 369584 149728 369636 149734
rect 369584 149670 369636 149676
rect 369688 7342 369716 172790
rect 369676 7336 369728 7342
rect 369676 7278 369728 7284
rect 369216 5160 369268 5166
rect 369216 5102 369268 5108
rect 368388 4548 368440 4554
rect 368388 4490 368440 4496
rect 367008 4480 367060 4486
rect 367008 4422 367060 4428
rect 368018 3496 368074 3505
rect 368018 3431 368074 3440
rect 368032 480 368060 3431
rect 369228 480 369256 5102
rect 369780 4622 369808 175100
rect 370240 172854 370268 175100
rect 370714 175086 371004 175114
rect 370228 172848 370280 172854
rect 370228 172790 370280 172796
rect 370976 148374 371004 175086
rect 371056 172848 371108 172854
rect 371056 172790 371108 172796
rect 370964 148368 371016 148374
rect 370964 148310 371016 148316
rect 370412 7948 370464 7954
rect 370412 7890 370464 7896
rect 369768 4616 369820 4622
rect 369768 4558 369820 4564
rect 370424 480 370452 7890
rect 371068 7410 371096 172790
rect 371056 7404 371108 7410
rect 371056 7346 371108 7352
rect 371160 4758 371188 175100
rect 371712 172854 371740 175100
rect 372186 175086 372476 175114
rect 371700 172848 371752 172854
rect 371700 172790 371752 172796
rect 372448 126274 372476 175086
rect 372632 172854 372660 175100
rect 372528 172848 372580 172854
rect 372528 172790 372580 172796
rect 372620 172848 372672 172854
rect 372620 172790 372672 172796
rect 372436 126268 372488 126274
rect 372436 126210 372488 126216
rect 372540 7478 372568 172790
rect 373092 172786 373120 175100
rect 373566 175086 373764 175114
rect 373080 172780 373132 172786
rect 373080 172722 373132 172728
rect 373736 146946 373764 175086
rect 374104 172922 374132 175100
rect 374092 172916 374144 172922
rect 374092 172858 374144 172864
rect 374564 172854 374592 175100
rect 375038 175086 375328 175114
rect 375196 172916 375248 172922
rect 375196 172858 375248 172864
rect 373908 172848 373960 172854
rect 373908 172790 373960 172796
rect 374552 172848 374604 172854
rect 374552 172790 374604 172796
rect 375104 172848 375156 172854
rect 375104 172790 375156 172796
rect 373816 172780 373868 172786
rect 373816 172722 373868 172728
rect 373724 146940 373776 146946
rect 373724 146882 373776 146888
rect 373828 7546 373856 172722
rect 373816 7540 373868 7546
rect 373816 7482 373868 7488
rect 372528 7472 372580 7478
rect 372528 7414 372580 7420
rect 372804 5092 372856 5098
rect 372804 5034 372856 5040
rect 371148 4752 371200 4758
rect 371148 4694 371200 4700
rect 371608 3596 371660 3602
rect 371608 3538 371660 3544
rect 371620 480 371648 3538
rect 372816 480 372844 5034
rect 373920 4690 373948 172790
rect 375116 8294 375144 172790
rect 375104 8288 375156 8294
rect 375104 8230 375156 8236
rect 374000 7880 374052 7886
rect 374000 7822 374052 7828
rect 373908 4684 373960 4690
rect 373908 4626 373960 4632
rect 374012 480 374040 7822
rect 375208 5506 375236 172858
rect 375196 5500 375248 5506
rect 375196 5442 375248 5448
rect 375300 3874 375328 175086
rect 375484 172922 375512 175100
rect 376050 175086 376340 175114
rect 376510 175086 376708 175114
rect 376312 173074 376340 175086
rect 376312 173046 376524 173074
rect 375472 172916 375524 172922
rect 375472 172858 375524 172864
rect 376496 8226 376524 173046
rect 376576 172916 376628 172922
rect 376576 172858 376628 172864
rect 376484 8220 376536 8226
rect 376484 8162 376536 8168
rect 376588 5438 376616 172858
rect 376576 5432 376628 5438
rect 376576 5374 376628 5380
rect 376392 5024 376444 5030
rect 376392 4966 376444 4972
rect 375288 3868 375340 3874
rect 375288 3810 375340 3816
rect 375194 3360 375250 3369
rect 375194 3295 375250 3304
rect 375208 480 375236 3295
rect 376404 480 376432 4966
rect 376680 3806 376708 175086
rect 376956 172922 376984 175100
rect 377784 173074 377812 175222
rect 377890 175086 378088 175114
rect 377784 173046 377904 173074
rect 376944 172916 376996 172922
rect 376944 172858 376996 172864
rect 377876 8158 377904 173046
rect 377956 172916 378008 172922
rect 377956 172858 378008 172864
rect 377864 8152 377916 8158
rect 377864 8094 377916 8100
rect 377588 7812 377640 7818
rect 377588 7754 377640 7760
rect 376668 3800 376720 3806
rect 376668 3742 376720 3748
rect 377600 480 377628 7754
rect 377968 5370 377996 172858
rect 377956 5364 378008 5370
rect 377956 5306 378008 5312
rect 378060 3738 378088 175086
rect 378428 172922 378456 175100
rect 378902 175086 379284 175114
rect 379362 175086 379468 175114
rect 378416 172916 378468 172922
rect 378416 172858 378468 172864
rect 378324 172780 378376 172786
rect 378324 172722 378376 172728
rect 378336 151842 378364 172722
rect 378140 151836 378192 151842
rect 378140 151778 378192 151784
rect 378324 151836 378376 151842
rect 378324 151778 378376 151784
rect 378152 151722 378180 151778
rect 378152 151694 378272 151722
rect 378244 142202 378272 151694
rect 378244 142174 378364 142202
rect 378336 132530 378364 142174
rect 378140 132524 378192 132530
rect 378140 132466 378192 132472
rect 378324 132524 378376 132530
rect 378324 132466 378376 132472
rect 378152 132410 378180 132466
rect 378152 132382 378272 132410
rect 378244 122890 378272 132382
rect 378244 122862 378364 122890
rect 378336 113218 378364 122862
rect 378140 113212 378192 113218
rect 378140 113154 378192 113160
rect 378324 113212 378376 113218
rect 378324 113154 378376 113160
rect 378152 113098 378180 113154
rect 378152 113070 378272 113098
rect 378244 103578 378272 113070
rect 378244 103550 378364 103578
rect 378336 93906 378364 103550
rect 378140 93900 378192 93906
rect 378140 93842 378192 93848
rect 378324 93900 378376 93906
rect 378324 93842 378376 93848
rect 378152 93786 378180 93842
rect 378152 93758 378272 93786
rect 378244 84266 378272 93758
rect 378244 84238 378364 84266
rect 378336 74594 378364 84238
rect 378140 74588 378192 74594
rect 378140 74530 378192 74536
rect 378324 74588 378376 74594
rect 378324 74530 378376 74536
rect 378152 74474 378180 74530
rect 378152 74446 378272 74474
rect 378244 64954 378272 74446
rect 378244 64926 378364 64954
rect 378336 55282 378364 64926
rect 378140 55276 378192 55282
rect 378140 55218 378192 55224
rect 378324 55276 378376 55282
rect 378324 55218 378376 55224
rect 378152 55162 378180 55218
rect 378152 55134 378272 55162
rect 378244 45642 378272 55134
rect 378244 45614 378364 45642
rect 378336 35970 378364 45614
rect 378140 35964 378192 35970
rect 378140 35906 378192 35912
rect 378324 35964 378376 35970
rect 378324 35906 378376 35912
rect 378152 26194 378180 35906
rect 378152 26166 378364 26194
rect 378336 16658 378364 26166
rect 378140 16652 378192 16658
rect 378140 16594 378192 16600
rect 378324 16652 378376 16658
rect 378324 16594 378376 16600
rect 378048 3732 378100 3738
rect 378048 3674 378100 3680
rect 378152 610 378180 16594
rect 379256 8090 379284 175086
rect 379336 172916 379388 172922
rect 379336 172858 379388 172864
rect 379244 8084 379296 8090
rect 379244 8026 379296 8032
rect 379348 5302 379376 172858
rect 379336 5296 379388 5302
rect 379336 5238 379388 5244
rect 379440 3670 379468 175086
rect 379808 172582 379836 175100
rect 380282 175086 380664 175114
rect 379796 172576 379848 172582
rect 379796 172518 379848 172524
rect 380636 8022 380664 175086
rect 380716 172576 380768 172582
rect 380716 172518 380768 172524
rect 380624 8016 380676 8022
rect 380624 7958 380676 7964
rect 380728 5234 380756 172518
rect 380716 5228 380768 5234
rect 380716 5170 380768 5176
rect 379980 4956 380032 4962
rect 379980 4898 380032 4904
rect 379428 3664 379480 3670
rect 379428 3606 379480 3612
rect 378140 604 378192 610
rect 378140 546 378192 552
rect 378784 604 378836 610
rect 378784 546 378836 552
rect 378796 480 378824 546
rect 379992 480 380020 4898
rect 380820 3602 380848 175100
rect 381280 172582 381308 175100
rect 381754 175086 382044 175114
rect 381268 172576 381320 172582
rect 381268 172518 381320 172524
rect 382016 7954 382044 175086
rect 382096 172576 382148 172582
rect 382096 172518 382148 172524
rect 382004 7948 382056 7954
rect 382004 7890 382056 7896
rect 381176 7744 381228 7750
rect 381176 7686 381228 7692
rect 380808 3596 380860 3602
rect 380808 3538 380860 3544
rect 381188 480 381216 7686
rect 382108 5166 382136 172518
rect 382096 5160 382148 5166
rect 382096 5102 382148 5108
rect 382200 3777 382228 175100
rect 382660 172582 382688 175100
rect 383226 175086 383516 175114
rect 382648 172576 382700 172582
rect 382648 172518 382700 172524
rect 383488 7886 383516 175086
rect 383672 172650 383700 175100
rect 383660 172644 383712 172650
rect 383660 172586 383712 172592
rect 384132 172582 384160 175100
rect 384606 175086 384804 175114
rect 383568 172576 383620 172582
rect 383568 172518 383620 172524
rect 384120 172576 384172 172582
rect 384120 172518 384172 172524
rect 383476 7880 383528 7886
rect 383476 7822 383528 7828
rect 383580 5098 383608 172518
rect 384776 7818 384804 175086
rect 385052 172650 385080 175100
rect 385408 172984 385460 172990
rect 385408 172926 385460 172932
rect 384948 172644 385000 172650
rect 384948 172586 385000 172592
rect 385040 172644 385092 172650
rect 385040 172586 385092 172592
rect 384856 172576 384908 172582
rect 384856 172518 384908 172524
rect 384764 7812 384816 7818
rect 384764 7754 384816 7760
rect 384672 7676 384724 7682
rect 384672 7618 384724 7624
rect 383568 5092 383620 5098
rect 383568 5034 383620 5040
rect 383568 4888 383620 4894
rect 383568 4830 383620 4836
rect 382186 3768 382242 3777
rect 382186 3703 382242 3712
rect 382372 3528 382424 3534
rect 382372 3470 382424 3476
rect 382384 480 382412 3470
rect 383580 480 383608 4830
rect 384684 480 384712 7618
rect 384868 5030 384896 172518
rect 384856 5024 384908 5030
rect 384856 4966 384908 4972
rect 384960 3534 384988 172586
rect 385420 166954 385448 172926
rect 385604 172582 385632 175100
rect 386078 175086 386184 175114
rect 385592 172576 385644 172582
rect 385592 172518 385644 172524
rect 385236 166926 385448 166954
rect 385236 164218 385264 166926
rect 385224 164212 385276 164218
rect 385224 164154 385276 164160
rect 385224 157344 385276 157350
rect 385224 157286 385276 157292
rect 385236 154578 385264 157286
rect 385236 154550 385356 154578
rect 385328 147694 385356 154550
rect 385132 147688 385184 147694
rect 385316 147688 385368 147694
rect 385184 147636 385264 147642
rect 385132 147630 385264 147636
rect 385316 147630 385368 147636
rect 385144 147614 385264 147630
rect 385236 144906 385264 147614
rect 385224 144900 385276 144906
rect 385224 144842 385276 144848
rect 385224 137964 385276 137970
rect 385224 137906 385276 137912
rect 385236 135266 385264 137906
rect 385236 135238 385356 135266
rect 385328 124234 385356 135238
rect 385040 124228 385092 124234
rect 385040 124170 385092 124176
rect 385316 124228 385368 124234
rect 385316 124170 385368 124176
rect 385052 119406 385080 124170
rect 385040 119400 385092 119406
rect 385040 119342 385092 119348
rect 385040 106344 385092 106350
rect 385040 106286 385092 106292
rect 385052 104854 385080 106286
rect 385040 104848 385092 104854
rect 385040 104790 385092 104796
rect 385132 93900 385184 93906
rect 385132 93842 385184 93848
rect 385144 84182 385172 93842
rect 385132 84176 385184 84182
rect 385132 84118 385184 84124
rect 385040 66292 385092 66298
rect 385040 66234 385092 66240
rect 385052 66201 385080 66234
rect 385038 66192 385094 66201
rect 385038 66127 385094 66136
rect 385130 60616 385186 60625
rect 385130 60551 385186 60560
rect 385144 51066 385172 60551
rect 385132 51060 385184 51066
rect 385132 51002 385184 51008
rect 385316 51060 385368 51066
rect 385316 51002 385368 51008
rect 385328 43466 385356 51002
rect 385328 43438 385448 43466
rect 385420 38622 385448 43438
rect 385408 38616 385460 38622
rect 385408 38558 385460 38564
rect 385316 29028 385368 29034
rect 385316 28970 385368 28976
rect 385328 22114 385356 28970
rect 385144 22086 385356 22114
rect 385144 19310 385172 22086
rect 385132 19304 385184 19310
rect 385132 19246 385184 19252
rect 385040 9716 385092 9722
rect 385040 9658 385092 9664
rect 385052 9602 385080 9658
rect 385052 9574 385172 9602
rect 384948 3528 385000 3534
rect 384948 3470 385000 3476
rect 385144 2650 385172 9574
rect 386156 7750 386184 175086
rect 386524 172650 386552 175100
rect 386328 172644 386380 172650
rect 386328 172586 386380 172592
rect 386512 172644 386564 172650
rect 386512 172586 386564 172592
rect 386236 172576 386288 172582
rect 386236 172518 386288 172524
rect 386144 7744 386196 7750
rect 386144 7686 386196 7692
rect 386248 4962 386276 172518
rect 386236 4956 386288 4962
rect 386236 4898 386288 4904
rect 386340 3641 386368 172586
rect 386984 172582 387012 175100
rect 387458 175086 387564 175114
rect 386972 172576 387024 172582
rect 386972 172518 387024 172524
rect 387536 7682 387564 175086
rect 387996 172650 388024 175100
rect 387708 172644 387760 172650
rect 387708 172586 387760 172592
rect 387984 172644 388036 172650
rect 387984 172586 388036 172592
rect 387616 172576 387668 172582
rect 387616 172518 387668 172524
rect 387524 7676 387576 7682
rect 387524 7618 387576 7624
rect 387628 4894 387656 172518
rect 387616 4888 387668 4894
rect 387616 4830 387668 4836
rect 387064 4820 387116 4826
rect 387064 4762 387116 4768
rect 386326 3632 386382 3641
rect 386326 3567 386382 3576
rect 385132 2644 385184 2650
rect 385132 2586 385184 2592
rect 385868 2644 385920 2650
rect 385868 2586 385920 2592
rect 385880 480 385908 2586
rect 387076 480 387104 4762
rect 387720 3505 387748 172586
rect 388456 172582 388484 175100
rect 388444 172576 388496 172582
rect 388444 172518 388496 172524
rect 388916 7614 388944 175100
rect 389376 172650 389404 175100
rect 389088 172644 389140 172650
rect 389088 172586 389140 172592
rect 389364 172644 389416 172650
rect 389364 172586 389416 172592
rect 390468 172644 390520 172650
rect 390468 172586 390520 172592
rect 388996 172576 389048 172582
rect 388996 172518 389048 172524
rect 388260 7608 388312 7614
rect 388260 7550 388312 7556
rect 388904 7608 388956 7614
rect 388904 7550 388956 7556
rect 387706 3496 387762 3505
rect 387706 3431 387762 3440
rect 388272 480 388300 7550
rect 389008 4826 389036 172518
rect 388996 4820 389048 4826
rect 388996 4762 389048 4768
rect 389100 3369 389128 172586
rect 390480 3466 390508 172586
rect 390560 170400 390612 170406
rect 390560 170342 390612 170348
rect 389456 3460 389508 3466
rect 389456 3402 389508 3408
rect 390468 3460 390520 3466
rect 390468 3402 390520 3408
rect 389086 3360 389142 3369
rect 389086 3295 389142 3304
rect 389468 480 389496 3402
rect 390572 626 390600 170342
rect 392596 30326 392624 182815
rect 392688 41410 392716 188119
rect 392780 77246 392808 198591
rect 392872 88330 392900 203895
rect 392964 124166 392992 214367
rect 393056 135250 393084 219671
rect 393148 158710 393176 224975
rect 393240 171086 393268 230143
rect 580172 229084 580224 229090
rect 580172 229026 580224 229032
rect 580184 228857 580212 229026
rect 580170 228848 580226 228857
rect 580170 228783 580226 228792
rect 580172 218000 580224 218006
rect 580172 217942 580224 217948
rect 580184 217025 580212 217942
rect 580170 217016 580226 217025
rect 580170 216951 580226 216960
rect 395344 208412 395396 208418
rect 395344 208354 395396 208360
rect 393962 193488 394018 193497
rect 393962 193423 394018 193432
rect 393228 171080 393280 171086
rect 393228 171022 393280 171028
rect 393136 158704 393188 158710
rect 393136 158646 393188 158652
rect 393320 156732 393372 156738
rect 393320 156674 393372 156680
rect 393044 135244 393096 135250
rect 393044 135186 393096 135192
rect 392952 124160 393004 124166
rect 392952 124102 393004 124108
rect 392860 88324 392912 88330
rect 392860 88266 392912 88272
rect 392768 77240 392820 77246
rect 392768 77182 392820 77188
rect 392676 41404 392728 41410
rect 392676 41346 392728 41352
rect 392584 30320 392636 30326
rect 392584 30262 392636 30268
rect 391848 7064 391900 7070
rect 391848 7006 391900 7012
rect 390572 598 390692 626
rect 390664 480 390692 598
rect 391860 480 391888 7006
rect 393332 3482 393360 156674
rect 393976 64870 394004 193423
rect 395356 111790 395384 208354
rect 579804 205624 579856 205630
rect 579804 205566 579856 205572
rect 579816 205329 579844 205566
rect 579802 205320 579858 205329
rect 579802 205255 579858 205264
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 519084 176724 519136 176730
rect 519084 176666 519136 176672
rect 409880 173868 409932 173874
rect 409880 173810 409932 173816
rect 402980 173120 403032 173126
rect 402980 173062 403032 173068
rect 396080 173052 396132 173058
rect 396080 172994 396132 173000
rect 395344 111784 395396 111790
rect 395344 111726 395396 111732
rect 393964 64864 394016 64870
rect 393964 64806 394016 64812
rect 395436 7132 395488 7138
rect 395436 7074 395488 7080
rect 393332 3454 394280 3482
rect 393044 2848 393096 2854
rect 393044 2790 393096 2796
rect 393056 480 393084 2790
rect 394252 480 394280 3454
rect 395448 480 395476 7074
rect 396092 3482 396120 172994
rect 397460 155304 397512 155310
rect 397460 155246 397512 155252
rect 397472 3482 397500 155246
rect 400312 153944 400364 153950
rect 400312 153886 400364 153892
rect 399024 8492 399076 8498
rect 399024 8434 399076 8440
rect 396092 3454 396672 3482
rect 397472 3454 397868 3482
rect 396644 480 396672 3454
rect 397840 480 397868 3454
rect 399036 480 399064 8434
rect 400324 3482 400352 153886
rect 402520 8560 402572 8566
rect 402520 8502 402572 8508
rect 400324 3454 401364 3482
rect 400220 2916 400272 2922
rect 400220 2858 400272 2864
rect 400232 480 400260 2858
rect 401336 480 401364 3454
rect 402532 480 402560 8502
rect 402992 3482 403020 173062
rect 404360 152584 404412 152590
rect 404360 152526 404412 152532
rect 404372 3482 404400 152526
rect 408500 151156 408552 151162
rect 408500 151098 408552 151104
rect 406108 8628 406160 8634
rect 406108 8570 406160 8576
rect 402992 3454 403756 3482
rect 404372 3454 404952 3482
rect 403728 480 403756 3454
rect 404924 480 404952 3454
rect 406120 480 406148 8570
rect 407304 2984 407356 2990
rect 407304 2926 407356 2932
rect 407316 480 407344 2926
rect 408512 480 408540 151098
rect 409696 8696 409748 8702
rect 409696 8638 409748 8644
rect 409708 480 409736 8638
rect 409892 3482 409920 173810
rect 416780 173800 416832 173806
rect 416780 173742 416832 173748
rect 411260 149796 411312 149802
rect 411260 149738 411312 149744
rect 411272 3482 411300 149738
rect 415400 148436 415452 148442
rect 415400 148378 415452 148384
rect 413284 8764 413336 8770
rect 413284 8706 413336 8712
rect 409892 3454 410932 3482
rect 411272 3454 412128 3482
rect 410904 480 410932 3454
rect 412100 480 412128 3454
rect 413296 480 413324 8706
rect 415412 3482 415440 148378
rect 415412 3454 415716 3482
rect 414480 3052 414532 3058
rect 414480 2994 414532 3000
rect 414492 480 414520 2994
rect 415688 480 415716 3454
rect 416792 3126 416820 173742
rect 425060 173732 425112 173738
rect 425060 173674 425112 173680
rect 418160 147008 418212 147014
rect 418160 146950 418212 146956
rect 416872 8832 416924 8838
rect 416872 8774 416924 8780
rect 416780 3120 416832 3126
rect 416780 3062 416832 3068
rect 416884 480 416912 8774
rect 418172 3482 418200 146950
rect 423956 9648 424008 9654
rect 423956 9590 424008 9596
rect 420368 8900 420420 8906
rect 420368 8842 420420 8848
rect 418172 3454 419212 3482
rect 417976 3120 418028 3126
rect 417976 3062 418028 3068
rect 417988 480 418016 3062
rect 419184 480 419212 3454
rect 420380 480 420408 8842
rect 422760 5636 422812 5642
rect 422760 5578 422812 5584
rect 421564 3052 421616 3058
rect 421564 2994 421616 3000
rect 421576 480 421604 2994
rect 422772 480 422800 5578
rect 423968 480 423996 9590
rect 425072 3482 425100 173674
rect 431960 173664 432012 173670
rect 431960 173606 432012 173612
rect 427544 9580 427596 9586
rect 427544 9522 427596 9528
rect 426348 5704 426400 5710
rect 426348 5646 426400 5652
rect 425072 3454 425192 3482
rect 425164 480 425192 3454
rect 426360 480 426388 5646
rect 427556 480 427584 9522
rect 431132 9512 431184 9518
rect 431132 9454 431184 9460
rect 429936 5772 429988 5778
rect 429936 5714 429988 5720
rect 428740 3188 428792 3194
rect 428740 3130 428792 3136
rect 428752 480 428780 3130
rect 429948 480 429976 5714
rect 431144 480 431172 9454
rect 431972 3482 432000 173606
rect 438860 173596 438912 173602
rect 438860 173538 438912 173544
rect 434628 9444 434680 9450
rect 434628 9386 434680 9392
rect 433524 5840 433576 5846
rect 433524 5782 433576 5788
rect 431972 3454 432368 3482
rect 432340 480 432368 3454
rect 433536 480 433564 5782
rect 434640 480 434668 9386
rect 438216 9376 438268 9382
rect 438216 9318 438268 9324
rect 437020 5908 437072 5914
rect 437020 5850 437072 5856
rect 435824 3256 435876 3262
rect 435824 3198 435876 3204
rect 435836 480 435864 3198
rect 437032 480 437060 5850
rect 438228 480 438256 9318
rect 438872 3482 438900 173538
rect 445760 173528 445812 173534
rect 445760 173470 445812 173476
rect 441804 9308 441856 9314
rect 441804 9250 441856 9256
rect 440608 5976 440660 5982
rect 440608 5918 440660 5924
rect 438872 3454 439452 3482
rect 439424 480 439452 3454
rect 440620 480 440648 5918
rect 441816 480 441844 9250
rect 445392 9240 445444 9246
rect 445392 9182 445444 9188
rect 444196 6044 444248 6050
rect 444196 5986 444248 5992
rect 443000 3324 443052 3330
rect 443000 3266 443052 3272
rect 443012 480 443040 3266
rect 444208 480 444236 5986
rect 445404 480 445432 9182
rect 445772 3482 445800 173470
rect 452660 173460 452712 173466
rect 452660 173402 452712 173408
rect 448980 9172 449032 9178
rect 448980 9114 449032 9120
rect 447784 6112 447836 6118
rect 447784 6054 447836 6060
rect 445772 3454 446628 3482
rect 446600 480 446628 3454
rect 447796 480 447824 6054
rect 448992 480 449020 9114
rect 452476 9104 452528 9110
rect 452476 9046 452528 9052
rect 451280 6860 451332 6866
rect 451280 6802 451332 6808
rect 450176 3392 450228 3398
rect 450176 3334 450228 3340
rect 450188 480 450216 3334
rect 451292 480 451320 6802
rect 452488 480 452516 9046
rect 452672 3482 452700 173402
rect 459560 173392 459612 173398
rect 459560 173334 459612 173340
rect 456064 9036 456116 9042
rect 456064 8978 456116 8984
rect 454868 6792 454920 6798
rect 454868 6734 454920 6740
rect 452672 3454 453712 3482
rect 453684 480 453712 3454
rect 454880 480 454908 6734
rect 456076 480 456104 8978
rect 458456 6724 458508 6730
rect 458456 6666 458508 6672
rect 457260 4140 457312 4146
rect 457260 4082 457312 4088
rect 457272 480 457300 4082
rect 458468 480 458496 6666
rect 459572 3398 459600 173334
rect 467840 173324 467892 173330
rect 467840 173266 467892 173272
rect 462320 137284 462372 137290
rect 462320 137226 462372 137232
rect 459652 8968 459704 8974
rect 459652 8910 459704 8916
rect 459560 3392 459612 3398
rect 459560 3334 459612 3340
rect 459664 480 459692 8910
rect 462044 6656 462096 6662
rect 462044 6598 462096 6604
rect 460848 3392 460900 3398
rect 460848 3334 460900 3340
rect 460860 480 460888 3334
rect 462056 480 462084 6598
rect 462332 3346 462360 137226
rect 466460 133204 466512 133210
rect 466460 133146 466512 133152
rect 465632 6588 465684 6594
rect 465632 6530 465684 6536
rect 464436 4072 464488 4078
rect 464436 4014 464488 4020
rect 462332 3318 463280 3346
rect 463252 480 463280 3318
rect 464448 480 464476 4014
rect 465644 480 465672 6530
rect 466472 3346 466500 133146
rect 467852 3482 467880 173266
rect 474740 173256 474792 173262
rect 474740 173198 474792 173204
rect 469220 135924 469272 135930
rect 469220 135866 469272 135872
rect 469128 6520 469180 6526
rect 469128 6462 469180 6468
rect 467852 3454 467972 3482
rect 466472 3318 466868 3346
rect 466840 480 466868 3318
rect 467944 480 467972 3454
rect 469140 480 469168 6462
rect 469232 3346 469260 135866
rect 473360 130416 473412 130422
rect 473360 130358 473412 130364
rect 472716 6452 472768 6458
rect 472716 6394 472768 6400
rect 471520 4004 471572 4010
rect 471520 3946 471572 3952
rect 469232 3318 470364 3346
rect 470336 480 470364 3318
rect 471532 480 471560 3946
rect 472728 480 472756 6394
rect 473372 3346 473400 130358
rect 474752 3346 474780 173198
rect 519096 173194 519124 176666
rect 481640 173188 481692 173194
rect 481640 173130 481692 173136
rect 519084 173188 519136 173194
rect 519084 173130 519136 173136
rect 580264 173188 580316 173194
rect 580264 173130 580316 173136
rect 477592 131776 477644 131782
rect 477592 131718 477644 131724
rect 476304 6384 476356 6390
rect 476304 6326 476356 6332
rect 473372 3318 473952 3346
rect 474752 3318 475148 3346
rect 473924 480 473952 3318
rect 475120 480 475148 3318
rect 476316 480 476344 6326
rect 477604 3482 477632 131718
rect 480260 127628 480312 127634
rect 480260 127570 480312 127576
rect 479892 6316 479944 6322
rect 479892 6258 479944 6264
rect 478696 3936 478748 3942
rect 478696 3878 478748 3884
rect 477512 3454 477632 3482
rect 477512 480 477540 3454
rect 478708 480 478736 3878
rect 479904 480 479932 6258
rect 480272 3346 480300 127570
rect 481652 3346 481680 173130
rect 483020 171828 483072 171834
rect 483020 171770 483072 171776
rect 483032 3346 483060 171770
rect 579896 171080 579948 171086
rect 579896 171022 579948 171028
rect 579908 170105 579936 171022
rect 579894 170096 579950 170105
rect 579894 170031 579950 170040
rect 485780 169040 485832 169046
rect 485780 168982 485832 168988
rect 484584 6248 484636 6254
rect 484584 6190 484636 6196
rect 480272 3318 481128 3346
rect 481652 3318 482324 3346
rect 483032 3318 483520 3346
rect 481100 480 481128 3318
rect 482296 480 482324 3318
rect 483492 480 483520 3318
rect 484596 480 484624 6190
rect 485792 3942 485820 168982
rect 489920 167680 489972 167686
rect 489920 167622 489972 167628
rect 485872 11756 485924 11762
rect 485872 11698 485924 11704
rect 485780 3936 485832 3942
rect 485780 3878 485832 3884
rect 485884 3482 485912 11698
rect 488540 10328 488592 10334
rect 488540 10270 488592 10276
rect 488172 6180 488224 6186
rect 488172 6122 488224 6128
rect 486976 3936 487028 3942
rect 486976 3878 487028 3884
rect 485792 3454 485912 3482
rect 485792 480 485820 3454
rect 486988 480 487016 3878
rect 488184 480 488212 6122
rect 488552 3346 488580 10270
rect 489932 3346 489960 167622
rect 494060 166320 494112 166326
rect 494060 166262 494112 166268
rect 491300 145580 491352 145586
rect 491300 145522 491352 145528
rect 491312 3346 491340 145522
rect 492680 129056 492732 129062
rect 492680 128998 492732 129004
rect 492692 3346 492720 128998
rect 494072 3482 494100 166262
rect 496820 164892 496872 164898
rect 496820 164834 496872 164840
rect 494152 14476 494204 14482
rect 494152 14418 494204 14424
rect 494164 3942 494192 14418
rect 495440 13116 495492 13122
rect 495440 13058 495492 13064
rect 494152 3936 494204 3942
rect 494152 3878 494204 3884
rect 495348 3936 495400 3942
rect 495348 3878 495400 3884
rect 494072 3454 494192 3482
rect 488552 3318 489408 3346
rect 489932 3318 490604 3346
rect 491312 3318 491800 3346
rect 492692 3318 492996 3346
rect 489380 480 489408 3318
rect 490576 480 490604 3318
rect 491772 480 491800 3318
rect 492968 480 492996 3318
rect 494164 480 494192 3454
rect 495360 480 495388 3878
rect 495452 3346 495480 13058
rect 496832 3346 496860 164834
rect 500960 163532 501012 163538
rect 500960 163474 501012 163480
rect 498200 141432 498252 141438
rect 498200 141374 498252 141380
rect 498212 3346 498240 141374
rect 499580 15904 499632 15910
rect 499580 15846 499632 15852
rect 499592 3346 499620 15846
rect 500972 3346 501000 163474
rect 503720 162172 503772 162178
rect 503720 162114 503772 162120
rect 502340 142860 502392 142866
rect 502340 142802 502392 142808
rect 502352 3482 502380 142802
rect 502432 17264 502484 17270
rect 502432 17206 502484 17212
rect 502444 3942 502472 17206
rect 502432 3936 502484 3942
rect 502432 3878 502484 3884
rect 503628 3936 503680 3942
rect 503628 3878 503680 3884
rect 502352 3454 502472 3482
rect 495452 3318 496584 3346
rect 496832 3318 497780 3346
rect 498212 3318 498976 3346
rect 499592 3318 500172 3346
rect 500972 3318 501276 3346
rect 496556 480 496584 3318
rect 497752 480 497780 3318
rect 498948 480 498976 3318
rect 500144 480 500172 3318
rect 501248 480 501276 3318
rect 502444 480 502472 3454
rect 503640 480 503668 3878
rect 503732 3346 503760 162114
rect 507860 160744 507912 160750
rect 507860 160686 507912 160692
rect 505100 144220 505152 144226
rect 505100 144162 505152 144168
rect 505112 3346 505140 144162
rect 506480 18624 506532 18630
rect 506480 18566 506532 18572
rect 506492 3346 506520 18566
rect 507872 3346 507900 160686
rect 512000 159384 512052 159390
rect 512000 159326 512052 159332
rect 509240 138712 509292 138718
rect 509240 138654 509292 138660
rect 509252 3482 509280 138654
rect 510620 19984 510672 19990
rect 510620 19926 510672 19932
rect 510632 3482 510660 19926
rect 509252 3454 509648 3482
rect 510632 3454 510844 3482
rect 503732 3318 504864 3346
rect 505112 3318 506060 3346
rect 506492 3318 507256 3346
rect 507872 3318 508452 3346
rect 504836 480 504864 3318
rect 506032 480 506060 3318
rect 507228 480 507256 3318
rect 508424 480 508452 3318
rect 509620 480 509648 3454
rect 510816 480 510844 3454
rect 512012 480 512040 159326
rect 580172 158704 580224 158710
rect 580172 158646 580224 158652
rect 580184 158409 580212 158646
rect 580170 158400 580226 158409
rect 580170 158335 580226 158344
rect 516140 156664 516192 156670
rect 516140 156606 516192 156612
rect 513380 153876 513432 153882
rect 513380 153818 513432 153824
rect 512092 140072 512144 140078
rect 512092 140014 512144 140020
rect 512104 3482 512132 140014
rect 513392 3482 513420 153818
rect 515588 4276 515640 4282
rect 515588 4218 515640 4224
rect 512104 3454 513236 3482
rect 513392 3454 514432 3482
rect 513208 480 513236 3454
rect 514404 480 514432 3454
rect 515600 480 515628 4218
rect 516152 3482 516180 156606
rect 520280 155236 520332 155242
rect 520280 155178 520332 155184
rect 517520 124908 517572 124914
rect 517520 124850 517572 124856
rect 517532 3482 517560 124850
rect 519084 4344 519136 4350
rect 519084 4286 519136 4292
rect 516152 3454 516824 3482
rect 517532 3454 517928 3482
rect 516796 480 516824 3454
rect 517900 480 517928 3454
rect 519096 480 519124 4286
rect 520292 480 520320 155178
rect 524420 152516 524472 152522
rect 524420 152458 524472 152464
rect 520372 21412 520424 21418
rect 520372 21354 520424 21360
rect 520384 610 520412 21354
rect 523868 7200 523920 7206
rect 523868 7142 523920 7148
rect 522672 4412 522724 4418
rect 522672 4354 522724 4360
rect 520372 604 520424 610
rect 520372 546 520424 552
rect 521476 604 521528 610
rect 521476 546 521528 552
rect 521488 480 521516 546
rect 522684 480 522712 4354
rect 523880 480 523908 7142
rect 524432 610 524460 152458
rect 528560 151088 528612 151094
rect 528560 151030 528612 151036
rect 527456 7268 527508 7274
rect 527456 7210 527508 7216
rect 526260 4480 526312 4486
rect 526260 4422 526312 4428
rect 524420 604 524472 610
rect 524420 546 524472 552
rect 525064 604 525116 610
rect 525064 546 525116 552
rect 525076 480 525104 546
rect 526272 480 526300 4422
rect 527468 480 527496 7210
rect 528572 592 528600 151030
rect 531320 149728 531372 149734
rect 531320 149670 531372 149676
rect 531044 7336 531096 7342
rect 531044 7278 531096 7284
rect 529848 4548 529900 4554
rect 529848 4490 529900 4496
rect 528572 564 528692 592
rect 528664 480 528692 564
rect 529860 480 529888 4490
rect 531056 480 531084 7278
rect 531332 610 531360 149670
rect 535460 148368 535512 148374
rect 535460 148310 535512 148316
rect 534540 7404 534592 7410
rect 534540 7346 534592 7352
rect 533436 4616 533488 4622
rect 533436 4558 533488 4564
rect 531320 604 531372 610
rect 531320 546 531372 552
rect 532240 604 532292 610
rect 532240 546 532292 552
rect 532252 480 532280 546
rect 533448 480 533476 4558
rect 534552 480 534580 7346
rect 535472 626 535500 148310
rect 542360 146940 542412 146946
rect 542360 146882 542412 146888
rect 538220 126268 538272 126274
rect 538220 126210 538272 126216
rect 538128 7472 538180 7478
rect 538128 7414 538180 7420
rect 536932 4752 536984 4758
rect 536932 4694 536984 4700
rect 535472 598 535684 626
rect 535656 592 535684 598
rect 535656 564 535776 592
rect 535748 480 535776 564
rect 536944 480 536972 4694
rect 538140 480 538168 7414
rect 538232 610 538260 126210
rect 541716 7540 541768 7546
rect 541716 7482 541768 7488
rect 540520 4684 540572 4690
rect 540520 4626 540572 4632
rect 538220 604 538272 610
rect 538220 546 538272 552
rect 539324 604 539376 610
rect 539324 546 539376 552
rect 539336 480 539364 546
rect 540532 480 540560 4626
rect 541728 480 541756 7482
rect 542372 610 542400 146882
rect 579896 135244 579948 135250
rect 579896 135186 579948 135192
rect 579908 134881 579936 135186
rect 579894 134872 579950 134881
rect 579894 134807 579950 134816
rect 579896 124160 579948 124166
rect 579896 124102 579948 124108
rect 579908 123185 579936 124102
rect 579894 123176 579950 123185
rect 579894 123111 579950 123120
rect 580172 111784 580224 111790
rect 580172 111726 580224 111732
rect 580184 111489 580212 111726
rect 580170 111480 580226 111489
rect 580170 111415 580226 111424
rect 579896 88324 579948 88330
rect 579896 88266 579948 88272
rect 579908 87961 579936 88266
rect 579894 87952 579950 87961
rect 579894 87887 579950 87896
rect 579896 77240 579948 77246
rect 579896 77182 579948 77188
rect 579908 76265 579936 77182
rect 579894 76256 579950 76265
rect 579894 76191 579950 76200
rect 580172 64864 580224 64870
rect 580172 64806 580224 64812
rect 580184 64569 580212 64806
rect 580170 64560 580226 64569
rect 580170 64495 580226 64504
rect 579896 41404 579948 41410
rect 579896 41346 579948 41352
rect 579908 41041 579936 41346
rect 579894 41032 579950 41041
rect 579894 40967 579950 40976
rect 579896 30320 579948 30326
rect 579896 30262 579948 30268
rect 579908 29345 579936 30262
rect 579894 29336 579950 29345
rect 579894 29271 579950 29280
rect 580276 17649 580304 173130
rect 580262 17640 580318 17649
rect 580262 17575 580318 17584
rect 545304 8288 545356 8294
rect 545304 8230 545356 8236
rect 544108 5500 544160 5506
rect 544108 5442 544160 5448
rect 542360 604 542412 610
rect 542360 546 542412 552
rect 542912 604 542964 610
rect 542912 546 542964 552
rect 542924 480 542952 546
rect 544120 480 544148 5442
rect 545316 480 545344 8230
rect 548892 8220 548944 8226
rect 548892 8162 548944 8168
rect 547696 5432 547748 5438
rect 547696 5374 547748 5380
rect 546500 3868 546552 3874
rect 546500 3810 546552 3816
rect 546512 480 546540 3810
rect 547708 480 547736 5374
rect 548904 480 548932 8162
rect 552388 8152 552440 8158
rect 552388 8094 552440 8100
rect 551192 5364 551244 5370
rect 551192 5306 551244 5312
rect 550088 3800 550140 3806
rect 550088 3742 550140 3748
rect 550100 480 550128 3742
rect 551204 480 551232 5306
rect 552400 480 552428 8094
rect 555976 8084 556028 8090
rect 555976 8026 556028 8032
rect 554780 5296 554832 5302
rect 554780 5238 554832 5244
rect 553584 3732 553636 3738
rect 553584 3674 553636 3680
rect 553596 480 553624 3674
rect 554792 480 554820 5238
rect 555988 480 556016 8026
rect 559564 8016 559616 8022
rect 559564 7958 559616 7964
rect 558368 5228 558420 5234
rect 558368 5170 558420 5176
rect 557172 3664 557224 3670
rect 557172 3606 557224 3612
rect 557184 480 557212 3606
rect 558380 480 558408 5170
rect 559576 480 559604 7958
rect 563152 7948 563204 7954
rect 563152 7890 563204 7896
rect 561956 5160 562008 5166
rect 561956 5102 562008 5108
rect 560760 3596 560812 3602
rect 560760 3538 560812 3544
rect 560772 480 560800 3538
rect 561968 480 561996 5102
rect 563164 480 563192 7890
rect 566740 7880 566792 7886
rect 566740 7822 566792 7828
rect 565544 5092 565596 5098
rect 565544 5034 565596 5040
rect 564346 3768 564402 3777
rect 564346 3703 564402 3712
rect 564360 480 564388 3703
rect 565556 480 565584 5034
rect 566752 480 566780 7822
rect 570236 7812 570288 7818
rect 570236 7754 570288 7760
rect 569040 5024 569092 5030
rect 569040 4966 569092 4972
rect 567844 3528 567896 3534
rect 567844 3470 567896 3476
rect 567856 480 567884 3470
rect 569052 480 569080 4966
rect 570248 480 570276 7754
rect 573824 7744 573876 7750
rect 573824 7686 573876 7692
rect 572628 4956 572680 4962
rect 572628 4898 572680 4904
rect 571430 3632 571486 3641
rect 571430 3567 571486 3576
rect 571444 480 571472 3567
rect 572640 480 572668 4898
rect 573836 480 573864 7686
rect 577412 7676 577464 7682
rect 577412 7618 577464 7624
rect 576216 4888 576268 4894
rect 576216 4830 576268 4836
rect 575018 3496 575074 3505
rect 575018 3431 575074 3440
rect 575032 480 575060 3431
rect 576228 480 576256 4830
rect 577424 480 577452 7618
rect 581000 7608 581052 7614
rect 581000 7550 581052 7556
rect 579804 4820 579856 4826
rect 579804 4762 579856 4768
rect 578606 3360 578662 3369
rect 578606 3295 578662 3304
rect 578620 480 578648 3295
rect 579816 480 579844 4762
rect 581012 480 581040 7550
rect 582196 3460 582248 3466
rect 582196 3402 582248 3408
rect 582208 480 582236 3402
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3330 682216 3386 682272
rect 3422 667936 3478 667992
rect 3054 624824 3110 624880
rect 3330 509904 3386 509960
rect 3330 452376 3386 452432
rect 3330 437960 3386 438016
rect 3330 423680 3386 423736
rect 3514 653520 3570 653576
rect 3606 610408 3662 610464
rect 3422 394984 3478 395040
rect 3698 595992 3754 596048
rect 4066 567296 4122 567352
rect 3790 553016 3846 553072
rect 3514 380568 3570 380624
rect 3882 538600 3938 538656
rect 3974 495488 4030 495544
rect 3606 366152 3662 366208
rect 4066 481072 4122 481128
rect 3698 337456 3754 337512
rect 3054 308760 3110 308816
rect 8114 531256 8170 531312
rect 8390 531256 8446 531312
rect 8114 511944 8170 512000
rect 8390 511944 8446 512000
rect 7930 473320 7986 473376
rect 8114 473320 8170 473376
rect 7838 415384 7894 415440
rect 8022 415384 8078 415440
rect 72974 608504 73030 608560
rect 73158 608504 73214 608560
rect 72698 531256 72754 531312
rect 72882 531256 72938 531312
rect 72606 511944 72662 512000
rect 72790 511944 72846 512000
rect 72882 434696 72938 434752
rect 73158 434696 73214 434752
rect 72882 425176 72938 425232
rect 72606 425040 72662 425096
rect 137834 531256 137890 531312
rect 138110 531256 138166 531312
rect 137834 511944 137890 512000
rect 138110 511944 138166 512000
rect 137650 482976 137706 483032
rect 137926 482976 137982 483032
rect 154210 482976 154266 483032
rect 154486 482976 154542 483032
rect 137374 454008 137430 454064
rect 137558 454008 137614 454064
rect 137558 415384 137614 415440
rect 137742 415384 137798 415440
rect 154118 415384 154174 415440
rect 154302 415384 154358 415440
rect 218886 695680 218942 695736
rect 219254 695544 219310 695600
rect 218978 540912 219034 540968
rect 219162 540912 219218 540968
rect 218978 531256 219034 531312
rect 219162 531256 219218 531312
rect 218886 511944 218942 512000
rect 219070 511944 219126 512000
rect 219162 434696 219218 434752
rect 219438 434696 219494 434752
rect 219162 425176 219218 425232
rect 218886 425040 218942 425096
rect 580170 697992 580226 698048
rect 391938 409128 391994 409184
rect 151818 408856 151874 408912
rect 392582 403824 392638 403880
rect 152370 403280 152426 403336
rect 391938 398520 391994 398576
rect 153106 397568 153162 397624
rect 391938 393352 391994 393408
rect 153106 391992 153162 392048
rect 391938 388048 391994 388104
rect 153106 386316 153108 386336
rect 153108 386316 153160 386336
rect 153160 386316 153162 386336
rect 153106 386280 153162 386316
rect 391938 382744 391994 382800
rect 152554 380704 152610 380760
rect 391938 377576 391994 377632
rect 152554 374992 152610 375048
rect 392674 372272 392730 372328
rect 152922 369416 152978 369472
rect 391938 367004 391940 367024
rect 391940 367004 391992 367024
rect 391992 367004 391994 367024
rect 391938 366968 391994 367004
rect 153106 363704 153162 363760
rect 391938 361800 391994 361856
rect 153106 358128 153162 358184
rect 391938 356496 391994 356552
rect 153106 352552 153162 352608
rect 391938 351192 391994 351248
rect 152922 346840 152978 346896
rect 391938 346024 391994 346080
rect 152554 341264 152610 341320
rect 153106 335552 153162 335608
rect 391938 335416 391994 335472
rect 391938 330112 391994 330168
rect 153106 329976 153162 330032
rect 391938 324944 391994 325000
rect 153106 324284 153162 324320
rect 153106 324264 153108 324284
rect 153108 324264 153160 324284
rect 153160 324264 153162 324284
rect 3790 323040 3846 323096
rect 391938 319640 391994 319696
rect 153106 318724 153108 318744
rect 153108 318724 153160 318744
rect 153160 318724 153162 318744
rect 153106 318688 153162 318724
rect 152370 312976 152426 313032
rect 391938 309168 391994 309224
rect 152554 307400 152610 307456
rect 391938 303864 391994 303920
rect 153106 301688 153162 301744
rect 392582 298560 392638 298616
rect 152738 296112 152794 296168
rect 3514 294344 3570 294400
rect 2962 280064 3018 280120
rect 392766 340720 392822 340776
rect 392674 293392 392730 293448
rect 152186 290536 152242 290592
rect 391938 288088 391994 288144
rect 152002 284824 152058 284880
rect 580170 686296 580226 686352
rect 580262 674600 580318 674656
rect 579894 639376 579950 639432
rect 392858 314336 392914 314392
rect 392766 282784 392822 282840
rect 152922 279248 152978 279304
rect 580170 592456 580226 592512
rect 580170 545536 580226 545592
rect 579986 498616 580042 498672
rect 579986 486784 580042 486840
rect 579986 463392 580042 463448
rect 579986 451696 580042 451752
rect 580170 439864 580226 439920
rect 580078 416472 580134 416528
rect 580078 404776 580134 404832
rect 580078 369552 580134 369608
rect 580078 357856 580134 357912
rect 580354 651072 580410 651128
rect 580446 627680 580502 627736
rect 580262 392944 580318 393000
rect 580170 322632 580226 322688
rect 579618 310800 579674 310856
rect 580538 604152 580594 604208
rect 580630 580760 580686 580816
rect 580722 557232 580778 557288
rect 580814 533840 580870 533896
rect 580906 510312 580962 510368
rect 580354 346024 580410 346080
rect 580262 299104 580318 299160
rect 392858 277616 392914 277672
rect 580170 275712 580226 275768
rect 152462 273536 152518 273592
rect 3422 265648 3478 265704
rect 3422 251232 3478 251288
rect 3146 208120 3202 208176
rect 3514 236952 3570 237008
rect 3514 222536 3570 222592
rect 3422 193840 3478 193896
rect 3054 179424 3110 179480
rect 3238 165008 3294 165064
rect 3330 136312 3386 136368
rect 3330 122032 3386 122088
rect 3054 78920 3110 78976
rect 3054 50088 3110 50144
rect 391938 272312 391994 272368
rect 153106 267960 153162 268016
rect 392582 267008 392638 267064
rect 579802 263880 579858 263936
rect 153106 262268 153162 262304
rect 153106 262248 153108 262268
rect 153108 262248 153160 262268
rect 153160 262248 153162 262268
rect 391938 261840 391994 261896
rect 152646 256672 152702 256728
rect 152554 245384 152610 245440
rect 152554 205944 152610 206000
rect 152002 200232 152058 200288
rect 152278 188944 152334 189000
rect 152462 183368 152518 183424
rect 3698 150728 3754 150784
rect 3606 107616 3662 107672
rect 3606 93200 3662 93256
rect 3514 64504 3570 64560
rect 3514 35844 3516 35864
rect 3516 35844 3568 35864
rect 3568 35844 3570 35864
rect 3514 35808 3570 35844
rect 3422 21392 3478 21448
rect 3422 7112 3478 7168
rect 5262 3304 5318 3360
rect 11242 3440 11298 3496
rect 19522 3576 19578 3632
rect 20718 3712 20774 3768
rect 391938 256536 391994 256592
rect 579802 252184 579858 252240
rect 392766 251232 392822 251288
rect 153106 250960 153162 251016
rect 392674 245928 392730 245984
rect 392582 240760 392638 240816
rect 152922 239672 152978 239728
rect 152738 222808 152794 222864
rect 152646 177792 152702 177848
rect 152830 194656 152886 194712
rect 392490 235456 392546 235512
rect 153106 234096 153162 234152
rect 153106 228520 153162 228576
rect 153014 217232 153070 217288
rect 153014 211520 153070 211576
rect 391938 209208 391994 209264
rect 393226 230152 393282 230208
rect 393134 224984 393190 225040
rect 393042 219680 393098 219736
rect 392950 214376 393006 214432
rect 392858 203904 392914 203960
rect 392766 198600 392822 198656
rect 392674 188128 392730 188184
rect 392582 182824 392638 182880
rect 391938 177656 391994 177712
rect 156418 3304 156474 3360
rect 157614 154536 157670 154592
rect 157798 154536 157854 154592
rect 157614 145016 157670 145072
rect 157614 144880 157670 144936
rect 158718 67632 158774 67688
rect 159086 164192 159142 164248
rect 159270 164192 159326 164248
rect 158994 145016 159050 145072
rect 158994 144880 159050 144936
rect 158994 67632 159050 67688
rect 158994 3440 159050 3496
rect 163042 143520 163098 143576
rect 163226 143540 163282 143576
rect 163226 143520 163228 143540
rect 163228 143520 163280 143540
rect 163280 143520 163282 143540
rect 162950 3712 163006 3768
rect 162858 3576 162914 3632
rect 168378 154536 168434 154592
rect 168378 133864 168434 133920
rect 168562 154536 168618 154592
rect 168562 133864 168618 133920
rect 172426 154536 172482 154592
rect 172610 154536 172666 154592
rect 179510 172488 179566 172544
rect 179694 172488 179750 172544
rect 179694 153176 179750 153232
rect 179878 153176 179934 153232
rect 183926 74704 183982 74760
rect 183834 74568 183890 74624
rect 185122 162832 185178 162888
rect 185306 162832 185362 162888
rect 193402 173848 193458 173904
rect 193678 173848 193734 173904
rect 193402 164192 193458 164248
rect 193586 164192 193642 164248
rect 193586 154672 193642 154728
rect 193494 154536 193550 154592
rect 194138 144744 194194 144800
rect 196254 135360 196310 135416
rect 196162 135224 196218 135280
rect 198738 154536 198794 154592
rect 198738 145016 198794 145072
rect 197634 135224 197690 135280
rect 197818 135224 197874 135280
rect 199014 154536 199070 154592
rect 200394 154672 200450 154728
rect 200394 154536 200450 154592
rect 206006 164212 206062 164248
rect 206006 164192 206008 164212
rect 206008 164192 206060 164212
rect 206060 164192 206062 164212
rect 206558 164192 206614 164248
rect 207202 154672 207258 154728
rect 207202 154556 207258 154592
rect 207202 154536 207204 154556
rect 207204 154536 207256 154556
rect 207256 154536 207258 154556
rect 207294 37440 207350 37496
rect 207386 37304 207442 37360
rect 209870 115912 209926 115968
rect 210146 115912 210202 115968
rect 209870 96600 209926 96656
rect 210146 96600 210202 96656
rect 217046 164212 217102 164248
rect 217046 164192 217048 164212
rect 217048 164192 217100 164212
rect 217100 164192 217102 164212
rect 217230 164192 217286 164248
rect 217046 145016 217102 145072
rect 217046 144880 217102 144936
rect 218242 125588 218298 125624
rect 218242 125568 218244 125588
rect 218244 125568 218296 125588
rect 218296 125568 218298 125588
rect 218426 125588 218482 125624
rect 218426 125568 218428 125588
rect 218428 125568 218480 125588
rect 218480 125568 218482 125588
rect 221094 162832 221150 162888
rect 221370 162832 221426 162888
rect 221002 125588 221058 125624
rect 221002 125568 221004 125588
rect 221004 125568 221056 125588
rect 221056 125568 221058 125588
rect 221186 125588 221242 125624
rect 221186 125568 221188 125588
rect 221188 125568 221240 125588
rect 221240 125568 221242 125588
rect 221094 113192 221150 113248
rect 221278 113192 221334 113248
rect 222566 164192 222622 164248
rect 222934 164192 222990 164248
rect 225234 143520 225290 143576
rect 225418 143520 225474 143576
rect 226706 164192 226762 164248
rect 227074 164192 227130 164248
rect 227994 164192 228050 164248
rect 228270 164192 228326 164248
rect 256514 57840 256570 57896
rect 256514 38528 256570 38584
rect 256790 154536 256846 154592
rect 256974 154556 257030 154592
rect 256974 154536 256976 154556
rect 256976 154536 257028 154556
rect 257028 154536 257030 154556
rect 256882 144880 256938 144936
rect 257158 144880 257214 144936
rect 256882 125568 256938 125624
rect 257158 125568 257214 125624
rect 256882 106256 256938 106312
rect 257158 106256 257214 106312
rect 256698 57840 256754 57896
rect 256698 38528 256754 38584
rect 299386 3712 299442 3768
rect 302146 3576 302202 3632
rect 303526 3440 303582 3496
rect 306286 3304 306342 3360
rect 357346 3712 357402 3768
rect 364522 3576 364578 3632
rect 368018 3440 368074 3496
rect 375194 3304 375250 3360
rect 382186 3712 382242 3768
rect 385038 66136 385094 66192
rect 385130 60560 385186 60616
rect 386326 3576 386382 3632
rect 387706 3440 387762 3496
rect 389086 3304 389142 3360
rect 580170 228792 580226 228848
rect 580170 216960 580226 217016
rect 393962 193432 394018 193488
rect 579802 205264 579858 205320
rect 580170 181872 580226 181928
rect 579894 170040 579950 170096
rect 580170 158344 580226 158400
rect 579894 134816 579950 134872
rect 579894 123120 579950 123176
rect 580170 111424 580226 111480
rect 579894 87896 579950 87952
rect 579894 76200 579950 76256
rect 580170 64504 580226 64560
rect 579894 40976 579950 41032
rect 579894 29280 579950 29336
rect 580262 17584 580318 17640
rect 564346 3712 564402 3768
rect 571430 3576 571486 3632
rect 575018 3440 575074 3496
rect 578606 3304 578662 3360
<< metal3 >>
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 218881 695738 218947 695741
rect 218881 695736 219450 695738
rect 218881 695680 218886 695736
rect 218942 695680 219450 695736
rect 218881 695678 219450 695680
rect 218881 695675 218947 695678
rect 219249 695602 219315 695605
rect 219390 695602 219450 695678
rect 219249 695600 219450 695602
rect 219249 695544 219254 695600
rect 219310 695544 219450 695600
rect 219249 695542 219450 695544
rect 219249 695539 219315 695542
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect -960 682274 480 682364
rect 3325 682274 3391 682277
rect -960 682272 3391 682274
rect -960 682216 3330 682272
rect 3386 682216 3391 682272
rect -960 682214 3391 682216
rect -960 682124 480 682214
rect 3325 682211 3391 682214
rect 580257 674658 580323 674661
rect 583520 674658 584960 674748
rect 580257 674656 584960 674658
rect 580257 674600 580262 674656
rect 580318 674600 584960 674656
rect 580257 674598 584960 674600
rect 580257 674595 580323 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3509 653578 3575 653581
rect -960 653576 3575 653578
rect -960 653520 3514 653576
rect 3570 653520 3575 653576
rect -960 653518 3575 653520
rect -960 653428 480 653518
rect 3509 653515 3575 653518
rect 580349 651130 580415 651133
rect 583520 651130 584960 651220
rect 580349 651128 584960 651130
rect 580349 651072 580354 651128
rect 580410 651072 584960 651128
rect 580349 651070 584960 651072
rect 580349 651067 580415 651070
rect 583520 650980 584960 651070
rect 579889 639434 579955 639437
rect 583520 639434 584960 639524
rect 579889 639432 584960 639434
rect 579889 639376 579894 639432
rect 579950 639376 584960 639432
rect 579889 639374 584960 639376
rect 579889 639371 579955 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 580441 627738 580507 627741
rect 583520 627738 584960 627828
rect 580441 627736 584960 627738
rect 580441 627680 580446 627736
rect 580502 627680 584960 627736
rect 580441 627678 584960 627680
rect 580441 627675 580507 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3049 624882 3115 624885
rect -960 624880 3115 624882
rect -960 624824 3054 624880
rect 3110 624824 3115 624880
rect -960 624822 3115 624824
rect -960 624732 480 624822
rect 3049 624819 3115 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3601 610466 3667 610469
rect -960 610464 3667 610466
rect -960 610408 3606 610464
rect 3662 610408 3667 610464
rect -960 610406 3667 610408
rect -960 610316 480 610406
rect 3601 610403 3667 610406
rect 72969 608562 73035 608565
rect 73153 608562 73219 608565
rect 72969 608560 73219 608562
rect 72969 608504 72974 608560
rect 73030 608504 73158 608560
rect 73214 608504 73219 608560
rect 72969 608502 73219 608504
rect 72969 608499 73035 608502
rect 73153 608499 73219 608502
rect 580533 604210 580599 604213
rect 583520 604210 584960 604300
rect 580533 604208 584960 604210
rect 580533 604152 580538 604208
rect 580594 604152 584960 604208
rect 580533 604150 584960 604152
rect 580533 604147 580599 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3693 596050 3759 596053
rect -960 596048 3759 596050
rect -960 595992 3698 596048
rect 3754 595992 3759 596048
rect -960 595990 3759 595992
rect -960 595900 480 595990
rect 3693 595987 3759 595990
rect 580165 592514 580231 592517
rect 583520 592514 584960 592604
rect 580165 592512 584960 592514
rect 580165 592456 580170 592512
rect 580226 592456 584960 592512
rect 580165 592454 584960 592456
rect 580165 592451 580231 592454
rect 583520 592364 584960 592454
rect -960 581620 480 581860
rect 580625 580818 580691 580821
rect 583520 580818 584960 580908
rect 580625 580816 584960 580818
rect 580625 580760 580630 580816
rect 580686 580760 584960 580816
rect 580625 580758 584960 580760
rect 580625 580755 580691 580758
rect 583520 580668 584960 580758
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 4061 567354 4127 567357
rect -960 567352 4127 567354
rect -960 567296 4066 567352
rect 4122 567296 4127 567352
rect -960 567294 4127 567296
rect -960 567204 480 567294
rect 4061 567291 4127 567294
rect 580717 557290 580783 557293
rect 583520 557290 584960 557380
rect 580717 557288 584960 557290
rect 580717 557232 580722 557288
rect 580778 557232 584960 557288
rect 580717 557230 584960 557232
rect 580717 557227 580783 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3785 553074 3851 553077
rect -960 553072 3851 553074
rect -960 553016 3790 553072
rect 3846 553016 3851 553072
rect -960 553014 3851 553016
rect -960 552924 480 553014
rect 3785 553011 3851 553014
rect 580165 545594 580231 545597
rect 583520 545594 584960 545684
rect 580165 545592 584960 545594
rect 580165 545536 580170 545592
rect 580226 545536 584960 545592
rect 580165 545534 584960 545536
rect 580165 545531 580231 545534
rect 583520 545444 584960 545534
rect 218973 540970 219039 540973
rect 219157 540970 219223 540973
rect 218973 540968 219223 540970
rect 218973 540912 218978 540968
rect 219034 540912 219162 540968
rect 219218 540912 219223 540968
rect 218973 540910 219223 540912
rect 218973 540907 219039 540910
rect 219157 540907 219223 540910
rect -960 538658 480 538748
rect 3877 538658 3943 538661
rect -960 538656 3943 538658
rect -960 538600 3882 538656
rect 3938 538600 3943 538656
rect -960 538598 3943 538600
rect -960 538508 480 538598
rect 3877 538595 3943 538598
rect 580809 533898 580875 533901
rect 583520 533898 584960 533988
rect 580809 533896 584960 533898
rect 580809 533840 580814 533896
rect 580870 533840 584960 533896
rect 580809 533838 584960 533840
rect 580809 533835 580875 533838
rect 583520 533748 584960 533838
rect 8109 531314 8175 531317
rect 8385 531314 8451 531317
rect 8109 531312 8451 531314
rect 8109 531256 8114 531312
rect 8170 531256 8390 531312
rect 8446 531256 8451 531312
rect 8109 531254 8451 531256
rect 8109 531251 8175 531254
rect 8385 531251 8451 531254
rect 72693 531314 72759 531317
rect 72877 531314 72943 531317
rect 72693 531312 72943 531314
rect 72693 531256 72698 531312
rect 72754 531256 72882 531312
rect 72938 531256 72943 531312
rect 72693 531254 72943 531256
rect 72693 531251 72759 531254
rect 72877 531251 72943 531254
rect 137829 531314 137895 531317
rect 138105 531314 138171 531317
rect 137829 531312 138171 531314
rect 137829 531256 137834 531312
rect 137890 531256 138110 531312
rect 138166 531256 138171 531312
rect 137829 531254 138171 531256
rect 137829 531251 137895 531254
rect 138105 531251 138171 531254
rect 218973 531314 219039 531317
rect 219157 531314 219223 531317
rect 218973 531312 219223 531314
rect 218973 531256 218978 531312
rect 219034 531256 219162 531312
rect 219218 531256 219223 531312
rect 218973 531254 219223 531256
rect 218973 531251 219039 531254
rect 219157 531251 219223 531254
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 8109 512002 8175 512005
rect 8385 512002 8451 512005
rect 8109 512000 8451 512002
rect 8109 511944 8114 512000
rect 8170 511944 8390 512000
rect 8446 511944 8451 512000
rect 8109 511942 8451 511944
rect 8109 511939 8175 511942
rect 8385 511939 8451 511942
rect 72601 512002 72667 512005
rect 72785 512002 72851 512005
rect 72601 512000 72851 512002
rect 72601 511944 72606 512000
rect 72662 511944 72790 512000
rect 72846 511944 72851 512000
rect 72601 511942 72851 511944
rect 72601 511939 72667 511942
rect 72785 511939 72851 511942
rect 137829 512002 137895 512005
rect 138105 512002 138171 512005
rect 137829 512000 138171 512002
rect 137829 511944 137834 512000
rect 137890 511944 138110 512000
rect 138166 511944 138171 512000
rect 137829 511942 138171 511944
rect 137829 511939 137895 511942
rect 138105 511939 138171 511942
rect 218881 512002 218947 512005
rect 219065 512002 219131 512005
rect 218881 512000 219131 512002
rect 218881 511944 218886 512000
rect 218942 511944 219070 512000
rect 219126 511944 219131 512000
rect 218881 511942 219131 511944
rect 218881 511939 218947 511942
rect 219065 511939 219131 511942
rect 580901 510370 580967 510373
rect 583520 510370 584960 510460
rect 580901 510368 584960 510370
rect 580901 510312 580906 510368
rect 580962 510312 584960 510368
rect 580901 510310 584960 510312
rect 580901 510307 580967 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3325 509962 3391 509965
rect -960 509960 3391 509962
rect -960 509904 3330 509960
rect 3386 509904 3391 509960
rect -960 509902 3391 509904
rect -960 509812 480 509902
rect 3325 509899 3391 509902
rect 579981 498674 580047 498677
rect 583520 498674 584960 498764
rect 579981 498672 584960 498674
rect 579981 498616 579986 498672
rect 580042 498616 584960 498672
rect 579981 498614 584960 498616
rect 579981 498611 580047 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 3969 495546 4035 495549
rect -960 495544 4035 495546
rect -960 495488 3974 495544
rect 4030 495488 4035 495544
rect -960 495486 4035 495488
rect -960 495396 480 495486
rect 3969 495483 4035 495486
rect 579981 486842 580047 486845
rect 583520 486842 584960 486932
rect 579981 486840 584960 486842
rect 579981 486784 579986 486840
rect 580042 486784 584960 486840
rect 579981 486782 584960 486784
rect 579981 486779 580047 486782
rect 583520 486692 584960 486782
rect 137645 483034 137711 483037
rect 137921 483034 137987 483037
rect 137645 483032 137987 483034
rect 137645 482976 137650 483032
rect 137706 482976 137926 483032
rect 137982 482976 137987 483032
rect 137645 482974 137987 482976
rect 137645 482971 137711 482974
rect 137921 482971 137987 482974
rect 154205 483034 154271 483037
rect 154481 483034 154547 483037
rect 154205 483032 154547 483034
rect 154205 482976 154210 483032
rect 154266 482976 154486 483032
rect 154542 482976 154547 483032
rect 154205 482974 154547 482976
rect 154205 482971 154271 482974
rect 154481 482971 154547 482974
rect -960 481130 480 481220
rect 4061 481130 4127 481133
rect -960 481128 4127 481130
rect -960 481072 4066 481128
rect 4122 481072 4127 481128
rect -960 481070 4127 481072
rect -960 480980 480 481070
rect 4061 481067 4127 481070
rect 583520 474996 584960 475236
rect 7925 473378 7991 473381
rect 8109 473378 8175 473381
rect 7925 473376 8175 473378
rect 7925 473320 7930 473376
rect 7986 473320 8114 473376
rect 8170 473320 8175 473376
rect 7925 473318 8175 473320
rect 7925 473315 7991 473318
rect 8109 473315 8175 473318
rect -960 466700 480 466940
rect 579981 463450 580047 463453
rect 583520 463450 584960 463540
rect 579981 463448 584960 463450
rect 579981 463392 579986 463448
rect 580042 463392 584960 463448
rect 579981 463390 584960 463392
rect 579981 463387 580047 463390
rect 583520 463300 584960 463390
rect 137369 454066 137435 454069
rect 137553 454066 137619 454069
rect 137369 454064 137619 454066
rect 137369 454008 137374 454064
rect 137430 454008 137558 454064
rect 137614 454008 137619 454064
rect 137369 454006 137619 454008
rect 137369 454003 137435 454006
rect 137553 454003 137619 454006
rect -960 452434 480 452524
rect 3325 452434 3391 452437
rect -960 452432 3391 452434
rect -960 452376 3330 452432
rect 3386 452376 3391 452432
rect -960 452374 3391 452376
rect -960 452284 480 452374
rect 3325 452371 3391 452374
rect 579981 451754 580047 451757
rect 583520 451754 584960 451844
rect 579981 451752 584960 451754
rect 579981 451696 579986 451752
rect 580042 451696 584960 451752
rect 579981 451694 584960 451696
rect 579981 451691 580047 451694
rect 583520 451604 584960 451694
rect 580165 439922 580231 439925
rect 583520 439922 584960 440012
rect 580165 439920 584960 439922
rect 580165 439864 580170 439920
rect 580226 439864 584960 439920
rect 580165 439862 584960 439864
rect 580165 439859 580231 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3325 438018 3391 438021
rect -960 438016 3391 438018
rect -960 437960 3330 438016
rect 3386 437960 3391 438016
rect -960 437958 3391 437960
rect -960 437868 480 437958
rect 3325 437955 3391 437958
rect 72877 434754 72943 434757
rect 73153 434754 73219 434757
rect 72877 434752 73219 434754
rect 72877 434696 72882 434752
rect 72938 434696 73158 434752
rect 73214 434696 73219 434752
rect 72877 434694 73219 434696
rect 72877 434691 72943 434694
rect 73153 434691 73219 434694
rect 219157 434754 219223 434757
rect 219433 434754 219499 434757
rect 219157 434752 219499 434754
rect 219157 434696 219162 434752
rect 219218 434696 219438 434752
rect 219494 434696 219499 434752
rect 219157 434694 219499 434696
rect 219157 434691 219223 434694
rect 219433 434691 219499 434694
rect 583520 428076 584960 428316
rect 72877 425234 72943 425237
rect 219157 425234 219223 425237
rect 72558 425232 72943 425234
rect 72558 425176 72882 425232
rect 72938 425176 72943 425232
rect 72558 425174 72943 425176
rect 72558 425101 72618 425174
rect 72877 425171 72943 425174
rect 218838 425232 219223 425234
rect 218838 425176 219162 425232
rect 219218 425176 219223 425232
rect 218838 425174 219223 425176
rect 218838 425101 218898 425174
rect 219157 425171 219223 425174
rect 72558 425096 72667 425101
rect 72558 425040 72606 425096
rect 72662 425040 72667 425096
rect 72558 425038 72667 425040
rect 218838 425096 218947 425101
rect 218838 425040 218886 425096
rect 218942 425040 218947 425096
rect 218838 425038 218947 425040
rect 72601 425035 72667 425038
rect 218881 425035 218947 425038
rect -960 423738 480 423828
rect 3325 423738 3391 423741
rect -960 423736 3391 423738
rect -960 423680 3330 423736
rect 3386 423680 3391 423736
rect -960 423678 3391 423680
rect -960 423588 480 423678
rect 3325 423675 3391 423678
rect 580073 416530 580139 416533
rect 583520 416530 584960 416620
rect 580073 416528 584960 416530
rect 580073 416472 580078 416528
rect 580134 416472 584960 416528
rect 580073 416470 584960 416472
rect 580073 416467 580139 416470
rect 583520 416380 584960 416470
rect 7833 415442 7899 415445
rect 8017 415442 8083 415445
rect 7833 415440 8083 415442
rect 7833 415384 7838 415440
rect 7894 415384 8022 415440
rect 8078 415384 8083 415440
rect 7833 415382 8083 415384
rect 7833 415379 7899 415382
rect 8017 415379 8083 415382
rect 137553 415442 137619 415445
rect 137737 415442 137803 415445
rect 137553 415440 137803 415442
rect 137553 415384 137558 415440
rect 137614 415384 137742 415440
rect 137798 415384 137803 415440
rect 137553 415382 137803 415384
rect 137553 415379 137619 415382
rect 137737 415379 137803 415382
rect 154113 415442 154179 415445
rect 154297 415442 154363 415445
rect 154113 415440 154363 415442
rect 154113 415384 154118 415440
rect 154174 415384 154302 415440
rect 154358 415384 154363 415440
rect 154113 415382 154363 415384
rect 154113 415379 154179 415382
rect 154297 415379 154363 415382
rect -960 409172 480 409412
rect 391933 409186 391999 409189
rect 389620 409184 391999 409186
rect 389620 409128 391938 409184
rect 391994 409128 391999 409184
rect 389620 409126 391999 409128
rect 391933 409123 391999 409126
rect 151813 408914 151879 408917
rect 151813 408912 155020 408914
rect 151813 408856 151818 408912
rect 151874 408856 155020 408912
rect 151813 408854 155020 408856
rect 151813 408851 151879 408854
rect 580073 404834 580139 404837
rect 583520 404834 584960 404924
rect 580073 404832 584960 404834
rect 580073 404776 580078 404832
rect 580134 404776 584960 404832
rect 580073 404774 584960 404776
rect 580073 404771 580139 404774
rect 583520 404684 584960 404774
rect 392577 403882 392643 403885
rect 389620 403880 392643 403882
rect 389620 403824 392582 403880
rect 392638 403824 392643 403880
rect 389620 403822 392643 403824
rect 392577 403819 392643 403822
rect 152365 403338 152431 403341
rect 152365 403336 155020 403338
rect 152365 403280 152370 403336
rect 152426 403280 155020 403336
rect 152365 403278 155020 403280
rect 152365 403275 152431 403278
rect 391933 398578 391999 398581
rect 389620 398576 391999 398578
rect 389620 398520 391938 398576
rect 391994 398520 391999 398576
rect 389620 398518 391999 398520
rect 391933 398515 391999 398518
rect 153101 397626 153167 397629
rect 153101 397624 155020 397626
rect 153101 397568 153106 397624
rect 153162 397568 155020 397624
rect 153101 397566 155020 397568
rect 153101 397563 153167 397566
rect -960 395042 480 395132
rect 3417 395042 3483 395045
rect -960 395040 3483 395042
rect -960 394984 3422 395040
rect 3478 394984 3483 395040
rect -960 394982 3483 394984
rect -960 394892 480 394982
rect 3417 394979 3483 394982
rect 391933 393410 391999 393413
rect 389620 393408 391999 393410
rect 389620 393352 391938 393408
rect 391994 393352 391999 393408
rect 389620 393350 391999 393352
rect 391933 393347 391999 393350
rect 580257 393002 580323 393005
rect 583520 393002 584960 393092
rect 580257 393000 584960 393002
rect 580257 392944 580262 393000
rect 580318 392944 584960 393000
rect 580257 392942 584960 392944
rect 580257 392939 580323 392942
rect 583520 392852 584960 392942
rect 153101 392050 153167 392053
rect 153101 392048 155020 392050
rect 153101 391992 153106 392048
rect 153162 391992 155020 392048
rect 153101 391990 155020 391992
rect 153101 391987 153167 391990
rect 391933 388106 391999 388109
rect 389620 388104 391999 388106
rect 389620 388048 391938 388104
rect 391994 388048 391999 388104
rect 389620 388046 391999 388048
rect 391933 388043 391999 388046
rect 153101 386338 153167 386341
rect 153101 386336 155020 386338
rect 153101 386280 153106 386336
rect 153162 386280 155020 386336
rect 153101 386278 155020 386280
rect 153101 386275 153167 386278
rect 391933 382802 391999 382805
rect 389620 382800 391999 382802
rect 389620 382744 391938 382800
rect 391994 382744 391999 382800
rect 389620 382742 391999 382744
rect 391933 382739 391999 382742
rect 583520 381156 584960 381396
rect 152549 380762 152615 380765
rect 152549 380760 155020 380762
rect -960 380626 480 380716
rect 152549 380704 152554 380760
rect 152610 380704 155020 380760
rect 152549 380702 155020 380704
rect 152549 380699 152615 380702
rect 3509 380626 3575 380629
rect -960 380624 3575 380626
rect -960 380568 3514 380624
rect 3570 380568 3575 380624
rect -960 380566 3575 380568
rect -960 380476 480 380566
rect 3509 380563 3575 380566
rect 391933 377634 391999 377637
rect 389620 377632 391999 377634
rect 389620 377576 391938 377632
rect 391994 377576 391999 377632
rect 389620 377574 391999 377576
rect 391933 377571 391999 377574
rect 152549 375050 152615 375053
rect 152549 375048 155020 375050
rect 152549 374992 152554 375048
rect 152610 374992 155020 375048
rect 152549 374990 155020 374992
rect 152549 374987 152615 374990
rect 392669 372330 392735 372333
rect 389620 372328 392735 372330
rect 389620 372272 392674 372328
rect 392730 372272 392735 372328
rect 389620 372270 392735 372272
rect 392669 372267 392735 372270
rect 580073 369610 580139 369613
rect 583520 369610 584960 369700
rect 580073 369608 584960 369610
rect 580073 369552 580078 369608
rect 580134 369552 584960 369608
rect 580073 369550 584960 369552
rect 580073 369547 580139 369550
rect 152917 369474 152983 369477
rect 152917 369472 155020 369474
rect 152917 369416 152922 369472
rect 152978 369416 155020 369472
rect 583520 369460 584960 369550
rect 152917 369414 155020 369416
rect 152917 369411 152983 369414
rect 391933 367026 391999 367029
rect 389620 367024 391999 367026
rect 389620 366968 391938 367024
rect 391994 366968 391999 367024
rect 389620 366966 391999 366968
rect 391933 366963 391999 366966
rect -960 366210 480 366300
rect 3601 366210 3667 366213
rect -960 366208 3667 366210
rect -960 366152 3606 366208
rect 3662 366152 3667 366208
rect -960 366150 3667 366152
rect -960 366060 480 366150
rect 3601 366147 3667 366150
rect 153101 363762 153167 363765
rect 153101 363760 155020 363762
rect 153101 363704 153106 363760
rect 153162 363704 155020 363760
rect 153101 363702 155020 363704
rect 153101 363699 153167 363702
rect 391933 361858 391999 361861
rect 389620 361856 391999 361858
rect 389620 361800 391938 361856
rect 391994 361800 391999 361856
rect 389620 361798 391999 361800
rect 391933 361795 391999 361798
rect 153101 358186 153167 358189
rect 153101 358184 155020 358186
rect 153101 358128 153106 358184
rect 153162 358128 155020 358184
rect 153101 358126 155020 358128
rect 153101 358123 153167 358126
rect 580073 357914 580139 357917
rect 583520 357914 584960 358004
rect 580073 357912 584960 357914
rect 580073 357856 580078 357912
rect 580134 357856 584960 357912
rect 580073 357854 584960 357856
rect 580073 357851 580139 357854
rect 583520 357764 584960 357854
rect 391933 356554 391999 356557
rect 389620 356552 391999 356554
rect 389620 356496 391938 356552
rect 391994 356496 391999 356552
rect 389620 356494 391999 356496
rect 391933 356491 391999 356494
rect 153101 352610 153167 352613
rect 153101 352608 155020 352610
rect 153101 352552 153106 352608
rect 153162 352552 155020 352608
rect 153101 352550 155020 352552
rect 153101 352547 153167 352550
rect -960 351780 480 352020
rect 391933 351250 391999 351253
rect 389620 351248 391999 351250
rect 389620 351192 391938 351248
rect 391994 351192 391999 351248
rect 389620 351190 391999 351192
rect 391933 351187 391999 351190
rect 152917 346898 152983 346901
rect 152917 346896 155020 346898
rect 152917 346840 152922 346896
rect 152978 346840 155020 346896
rect 152917 346838 155020 346840
rect 152917 346835 152983 346838
rect 391933 346082 391999 346085
rect 389620 346080 391999 346082
rect 389620 346024 391938 346080
rect 391994 346024 391999 346080
rect 389620 346022 391999 346024
rect 391933 346019 391999 346022
rect 580349 346082 580415 346085
rect 583520 346082 584960 346172
rect 580349 346080 584960 346082
rect 580349 346024 580354 346080
rect 580410 346024 584960 346080
rect 580349 346022 584960 346024
rect 580349 346019 580415 346022
rect 583520 345932 584960 346022
rect 152549 341322 152615 341325
rect 152549 341320 155020 341322
rect 152549 341264 152554 341320
rect 152610 341264 155020 341320
rect 152549 341262 155020 341264
rect 152549 341259 152615 341262
rect 392761 340778 392827 340781
rect 389620 340776 392827 340778
rect 389620 340720 392766 340776
rect 392822 340720 392827 340776
rect 389620 340718 392827 340720
rect 392761 340715 392827 340718
rect -960 337514 480 337604
rect 3693 337514 3759 337517
rect -960 337512 3759 337514
rect -960 337456 3698 337512
rect 3754 337456 3759 337512
rect -960 337454 3759 337456
rect -960 337364 480 337454
rect 3693 337451 3759 337454
rect 153101 335610 153167 335613
rect 153101 335608 155020 335610
rect 153101 335552 153106 335608
rect 153162 335552 155020 335608
rect 153101 335550 155020 335552
rect 153101 335547 153167 335550
rect 391933 335474 391999 335477
rect 389620 335472 391999 335474
rect 389620 335416 391938 335472
rect 391994 335416 391999 335472
rect 389620 335414 391999 335416
rect 391933 335411 391999 335414
rect 583520 334236 584960 334476
rect 391933 330170 391999 330173
rect 389620 330168 391999 330170
rect 389620 330112 391938 330168
rect 391994 330112 391999 330168
rect 389620 330110 391999 330112
rect 391933 330107 391999 330110
rect 153101 330034 153167 330037
rect 153101 330032 155020 330034
rect 153101 329976 153106 330032
rect 153162 329976 155020 330032
rect 153101 329974 155020 329976
rect 153101 329971 153167 329974
rect 391933 325002 391999 325005
rect 389620 325000 391999 325002
rect 389620 324944 391938 325000
rect 391994 324944 391999 325000
rect 389620 324942 391999 324944
rect 391933 324939 391999 324942
rect 153101 324322 153167 324325
rect 153101 324320 155020 324322
rect 153101 324264 153106 324320
rect 153162 324264 155020 324320
rect 153101 324262 155020 324264
rect 153101 324259 153167 324262
rect -960 323098 480 323188
rect 3785 323098 3851 323101
rect -960 323096 3851 323098
rect -960 323040 3790 323096
rect 3846 323040 3851 323096
rect -960 323038 3851 323040
rect -960 322948 480 323038
rect 3785 323035 3851 323038
rect 580165 322690 580231 322693
rect 583520 322690 584960 322780
rect 580165 322688 584960 322690
rect 580165 322632 580170 322688
rect 580226 322632 584960 322688
rect 580165 322630 584960 322632
rect 580165 322627 580231 322630
rect 583520 322540 584960 322630
rect 391933 319698 391999 319701
rect 389620 319696 391999 319698
rect 389620 319640 391938 319696
rect 391994 319640 391999 319696
rect 389620 319638 391999 319640
rect 391933 319635 391999 319638
rect 153101 318746 153167 318749
rect 153101 318744 155020 318746
rect 153101 318688 153106 318744
rect 153162 318688 155020 318744
rect 153101 318686 155020 318688
rect 153101 318683 153167 318686
rect 392853 314394 392919 314397
rect 389620 314392 392919 314394
rect 389620 314336 392858 314392
rect 392914 314336 392919 314392
rect 389620 314334 392919 314336
rect 392853 314331 392919 314334
rect 152365 313034 152431 313037
rect 152365 313032 155020 313034
rect 152365 312976 152370 313032
rect 152426 312976 155020 313032
rect 152365 312974 155020 312976
rect 152365 312971 152431 312974
rect 579613 310858 579679 310861
rect 583520 310858 584960 310948
rect 579613 310856 584960 310858
rect 579613 310800 579618 310856
rect 579674 310800 584960 310856
rect 579613 310798 584960 310800
rect 579613 310795 579679 310798
rect 583520 310708 584960 310798
rect 391933 309226 391999 309229
rect 389620 309224 391999 309226
rect 389620 309168 391938 309224
rect 391994 309168 391999 309224
rect 389620 309166 391999 309168
rect 391933 309163 391999 309166
rect -960 308818 480 308908
rect 3049 308818 3115 308821
rect -960 308816 3115 308818
rect -960 308760 3054 308816
rect 3110 308760 3115 308816
rect -960 308758 3115 308760
rect -960 308668 480 308758
rect 3049 308755 3115 308758
rect 152549 307458 152615 307461
rect 152549 307456 155020 307458
rect 152549 307400 152554 307456
rect 152610 307400 155020 307456
rect 152549 307398 155020 307400
rect 152549 307395 152615 307398
rect 391933 303922 391999 303925
rect 389620 303920 391999 303922
rect 389620 303864 391938 303920
rect 391994 303864 391999 303920
rect 389620 303862 391999 303864
rect 391933 303859 391999 303862
rect 153101 301746 153167 301749
rect 153101 301744 155020 301746
rect 153101 301688 153106 301744
rect 153162 301688 155020 301744
rect 153101 301686 155020 301688
rect 153101 301683 153167 301686
rect 580257 299162 580323 299165
rect 583520 299162 584960 299252
rect 580257 299160 584960 299162
rect 580257 299104 580262 299160
rect 580318 299104 584960 299160
rect 580257 299102 584960 299104
rect 580257 299099 580323 299102
rect 583520 299012 584960 299102
rect 392577 298618 392643 298621
rect 389620 298616 392643 298618
rect 389620 298560 392582 298616
rect 392638 298560 392643 298616
rect 389620 298558 392643 298560
rect 392577 298555 392643 298558
rect 152733 296170 152799 296173
rect 152733 296168 155020 296170
rect 152733 296112 152738 296168
rect 152794 296112 155020 296168
rect 152733 296110 155020 296112
rect 152733 296107 152799 296110
rect -960 294402 480 294492
rect 3509 294402 3575 294405
rect -960 294400 3575 294402
rect -960 294344 3514 294400
rect 3570 294344 3575 294400
rect -960 294342 3575 294344
rect -960 294252 480 294342
rect 3509 294339 3575 294342
rect 392669 293450 392735 293453
rect 389620 293448 392735 293450
rect 389620 293392 392674 293448
rect 392730 293392 392735 293448
rect 389620 293390 392735 293392
rect 392669 293387 392735 293390
rect 152181 290594 152247 290597
rect 152181 290592 155020 290594
rect 152181 290536 152186 290592
rect 152242 290536 155020 290592
rect 152181 290534 155020 290536
rect 152181 290531 152247 290534
rect 391933 288146 391999 288149
rect 389620 288144 391999 288146
rect 389620 288088 391938 288144
rect 391994 288088 391999 288144
rect 389620 288086 391999 288088
rect 391933 288083 391999 288086
rect 583520 287316 584960 287556
rect 151997 284882 152063 284885
rect 151997 284880 155020 284882
rect 151997 284824 152002 284880
rect 152058 284824 155020 284880
rect 151997 284822 155020 284824
rect 151997 284819 152063 284822
rect 392761 282842 392827 282845
rect 389620 282840 392827 282842
rect 389620 282784 392766 282840
rect 392822 282784 392827 282840
rect 389620 282782 392827 282784
rect 392761 282779 392827 282782
rect -960 280122 480 280212
rect 2957 280122 3023 280125
rect -960 280120 3023 280122
rect -960 280064 2962 280120
rect 3018 280064 3023 280120
rect -960 280062 3023 280064
rect -960 279972 480 280062
rect 2957 280059 3023 280062
rect 152917 279306 152983 279309
rect 152917 279304 155020 279306
rect 152917 279248 152922 279304
rect 152978 279248 155020 279304
rect 152917 279246 155020 279248
rect 152917 279243 152983 279246
rect 392853 277674 392919 277677
rect 389620 277672 392919 277674
rect 389620 277616 392858 277672
rect 392914 277616 392919 277672
rect 389620 277614 392919 277616
rect 392853 277611 392919 277614
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 152457 273594 152523 273597
rect 152457 273592 155020 273594
rect 152457 273536 152462 273592
rect 152518 273536 155020 273592
rect 152457 273534 155020 273536
rect 152457 273531 152523 273534
rect 391933 272370 391999 272373
rect 389620 272368 391999 272370
rect 389620 272312 391938 272368
rect 391994 272312 391999 272368
rect 389620 272310 391999 272312
rect 391933 272307 391999 272310
rect 153101 268018 153167 268021
rect 153101 268016 155020 268018
rect 153101 267960 153106 268016
rect 153162 267960 155020 268016
rect 153101 267958 155020 267960
rect 153101 267955 153167 267958
rect 392577 267066 392643 267069
rect 389620 267064 392643 267066
rect 389620 267008 392582 267064
rect 392638 267008 392643 267064
rect 389620 267006 392643 267008
rect 392577 267003 392643 267006
rect -960 265706 480 265796
rect 3417 265706 3483 265709
rect -960 265704 3483 265706
rect -960 265648 3422 265704
rect 3478 265648 3483 265704
rect -960 265646 3483 265648
rect -960 265556 480 265646
rect 3417 265643 3483 265646
rect 579797 263938 579863 263941
rect 583520 263938 584960 264028
rect 579797 263936 584960 263938
rect 579797 263880 579802 263936
rect 579858 263880 584960 263936
rect 579797 263878 584960 263880
rect 579797 263875 579863 263878
rect 583520 263788 584960 263878
rect 153101 262306 153167 262309
rect 153101 262304 155020 262306
rect 153101 262248 153106 262304
rect 153162 262248 155020 262304
rect 153101 262246 155020 262248
rect 153101 262243 153167 262246
rect 391933 261898 391999 261901
rect 389620 261896 391999 261898
rect 389620 261840 391938 261896
rect 391994 261840 391999 261896
rect 389620 261838 391999 261840
rect 391933 261835 391999 261838
rect 152641 256730 152707 256733
rect 152641 256728 155020 256730
rect 152641 256672 152646 256728
rect 152702 256672 155020 256728
rect 152641 256670 155020 256672
rect 152641 256667 152707 256670
rect 391933 256594 391999 256597
rect 389620 256592 391999 256594
rect 389620 256536 391938 256592
rect 391994 256536 391999 256592
rect 389620 256534 391999 256536
rect 391933 256531 391999 256534
rect 579797 252242 579863 252245
rect 583520 252242 584960 252332
rect 579797 252240 584960 252242
rect 579797 252184 579802 252240
rect 579858 252184 584960 252240
rect 579797 252182 584960 252184
rect 579797 252179 579863 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3417 251290 3483 251293
rect 392761 251290 392827 251293
rect -960 251288 3483 251290
rect -960 251232 3422 251288
rect 3478 251232 3483 251288
rect -960 251230 3483 251232
rect 389620 251288 392827 251290
rect 389620 251232 392766 251288
rect 392822 251232 392827 251288
rect 389620 251230 392827 251232
rect -960 251140 480 251230
rect 3417 251227 3483 251230
rect 392761 251227 392827 251230
rect 153101 251018 153167 251021
rect 153101 251016 155020 251018
rect 153101 250960 153106 251016
rect 153162 250960 155020 251016
rect 153101 250958 155020 250960
rect 153101 250955 153167 250958
rect 392669 245986 392735 245989
rect 389620 245984 392735 245986
rect 389620 245928 392674 245984
rect 392730 245928 392735 245984
rect 389620 245926 392735 245928
rect 392669 245923 392735 245926
rect 152549 245442 152615 245445
rect 152549 245440 155020 245442
rect 152549 245384 152554 245440
rect 152610 245384 155020 245440
rect 152549 245382 155020 245384
rect 152549 245379 152615 245382
rect 392577 240818 392643 240821
rect 389620 240816 392643 240818
rect 389620 240760 392582 240816
rect 392638 240760 392643 240816
rect 389620 240758 392643 240760
rect 392577 240755 392643 240758
rect 583520 240396 584960 240636
rect 152917 239730 152983 239733
rect 152917 239728 155020 239730
rect 152917 239672 152922 239728
rect 152978 239672 155020 239728
rect 152917 239670 155020 239672
rect 152917 239667 152983 239670
rect -960 237010 480 237100
rect 3509 237010 3575 237013
rect -960 237008 3575 237010
rect -960 236952 3514 237008
rect 3570 236952 3575 237008
rect -960 236950 3575 236952
rect -960 236860 480 236950
rect 3509 236947 3575 236950
rect 392485 235514 392551 235517
rect 389620 235512 392551 235514
rect 389620 235456 392490 235512
rect 392546 235456 392551 235512
rect 389620 235454 392551 235456
rect 392485 235451 392551 235454
rect 153101 234154 153167 234157
rect 153101 234152 155020 234154
rect 153101 234096 153106 234152
rect 153162 234096 155020 234152
rect 153101 234094 155020 234096
rect 153101 234091 153167 234094
rect 393221 230210 393287 230213
rect 389620 230208 393287 230210
rect 389620 230152 393226 230208
rect 393282 230152 393287 230208
rect 389620 230150 393287 230152
rect 393221 230147 393287 230150
rect 580165 228850 580231 228853
rect 583520 228850 584960 228940
rect 580165 228848 584960 228850
rect 580165 228792 580170 228848
rect 580226 228792 584960 228848
rect 580165 228790 584960 228792
rect 580165 228787 580231 228790
rect 583520 228700 584960 228790
rect 153101 228578 153167 228581
rect 153101 228576 155020 228578
rect 153101 228520 153106 228576
rect 153162 228520 155020 228576
rect 153101 228518 155020 228520
rect 153101 228515 153167 228518
rect 393129 225042 393195 225045
rect 389620 225040 393195 225042
rect 389620 224984 393134 225040
rect 393190 224984 393195 225040
rect 389620 224982 393195 224984
rect 393129 224979 393195 224982
rect 152733 222866 152799 222869
rect 152733 222864 155020 222866
rect 152733 222808 152738 222864
rect 152794 222808 155020 222864
rect 152733 222806 155020 222808
rect 152733 222803 152799 222806
rect -960 222594 480 222684
rect 3509 222594 3575 222597
rect -960 222592 3575 222594
rect -960 222536 3514 222592
rect 3570 222536 3575 222592
rect -960 222534 3575 222536
rect -960 222444 480 222534
rect 3509 222531 3575 222534
rect 393037 219738 393103 219741
rect 389620 219736 393103 219738
rect 389620 219680 393042 219736
rect 393098 219680 393103 219736
rect 389620 219678 393103 219680
rect 393037 219675 393103 219678
rect 153009 217290 153075 217293
rect 153009 217288 155020 217290
rect 153009 217232 153014 217288
rect 153070 217232 155020 217288
rect 153009 217230 155020 217232
rect 153009 217227 153075 217230
rect 580165 217018 580231 217021
rect 583520 217018 584960 217108
rect 580165 217016 584960 217018
rect 580165 216960 580170 217016
rect 580226 216960 584960 217016
rect 580165 216958 584960 216960
rect 580165 216955 580231 216958
rect 583520 216868 584960 216958
rect 392945 214434 393011 214437
rect 389620 214432 393011 214434
rect 389620 214376 392950 214432
rect 393006 214376 393011 214432
rect 389620 214374 393011 214376
rect 392945 214371 393011 214374
rect 153009 211578 153075 211581
rect 153009 211576 155020 211578
rect 153009 211520 153014 211576
rect 153070 211520 155020 211576
rect 153009 211518 155020 211520
rect 153009 211515 153075 211518
rect 391933 209266 391999 209269
rect 389620 209264 391999 209266
rect 389620 209208 391938 209264
rect 391994 209208 391999 209264
rect 389620 209206 391999 209208
rect 391933 209203 391999 209206
rect -960 208178 480 208268
rect 3141 208178 3207 208181
rect -960 208176 3207 208178
rect -960 208120 3146 208176
rect 3202 208120 3207 208176
rect -960 208118 3207 208120
rect -960 208028 480 208118
rect 3141 208115 3207 208118
rect 152549 206002 152615 206005
rect 152549 206000 155020 206002
rect 152549 205944 152554 206000
rect 152610 205944 155020 206000
rect 152549 205942 155020 205944
rect 152549 205939 152615 205942
rect 579797 205322 579863 205325
rect 583520 205322 584960 205412
rect 579797 205320 584960 205322
rect 579797 205264 579802 205320
rect 579858 205264 584960 205320
rect 579797 205262 584960 205264
rect 579797 205259 579863 205262
rect 583520 205172 584960 205262
rect 392853 203962 392919 203965
rect 389620 203960 392919 203962
rect 389620 203904 392858 203960
rect 392914 203904 392919 203960
rect 389620 203902 392919 203904
rect 392853 203899 392919 203902
rect 151997 200290 152063 200293
rect 151997 200288 155020 200290
rect 151997 200232 152002 200288
rect 152058 200232 155020 200288
rect 151997 200230 155020 200232
rect 151997 200227 152063 200230
rect 392761 198658 392827 198661
rect 389620 198656 392827 198658
rect 389620 198600 392766 198656
rect 392822 198600 392827 198656
rect 389620 198598 392827 198600
rect 392761 198595 392827 198598
rect 152825 194714 152891 194717
rect 152825 194712 155020 194714
rect 152825 194656 152830 194712
rect 152886 194656 155020 194712
rect 152825 194654 155020 194656
rect 152825 194651 152891 194654
rect -960 193898 480 193988
rect 3417 193898 3483 193901
rect -960 193896 3483 193898
rect -960 193840 3422 193896
rect 3478 193840 3483 193896
rect -960 193838 3483 193840
rect -960 193748 480 193838
rect 3417 193835 3483 193838
rect 393957 193490 394023 193493
rect 389620 193488 394023 193490
rect 389620 193432 393962 193488
rect 394018 193432 394023 193488
rect 583520 193476 584960 193716
rect 389620 193430 394023 193432
rect 393957 193427 394023 193430
rect 152273 189002 152339 189005
rect 152273 189000 155020 189002
rect 152273 188944 152278 189000
rect 152334 188944 155020 189000
rect 152273 188942 155020 188944
rect 152273 188939 152339 188942
rect 392669 188186 392735 188189
rect 389620 188184 392735 188186
rect 389620 188128 392674 188184
rect 392730 188128 392735 188184
rect 389620 188126 392735 188128
rect 392669 188123 392735 188126
rect 152457 183426 152523 183429
rect 152457 183424 155020 183426
rect 152457 183368 152462 183424
rect 152518 183368 155020 183424
rect 152457 183366 155020 183368
rect 152457 183363 152523 183366
rect 392577 182882 392643 182885
rect 389620 182880 392643 182882
rect 389620 182824 392582 182880
rect 392638 182824 392643 182880
rect 389620 182822 392643 182824
rect 392577 182819 392643 182822
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 3049 179482 3115 179485
rect -960 179480 3115 179482
rect -960 179424 3054 179480
rect 3110 179424 3115 179480
rect -960 179422 3115 179424
rect -960 179332 480 179422
rect 3049 179419 3115 179422
rect 152641 177850 152707 177853
rect 152641 177848 155020 177850
rect 152641 177792 152646 177848
rect 152702 177792 155020 177848
rect 152641 177790 155020 177792
rect 152641 177787 152707 177790
rect 391933 177714 391999 177717
rect 389620 177712 391999 177714
rect 389620 177656 391938 177712
rect 391994 177656 391999 177712
rect 389620 177654 391999 177656
rect 391933 177651 391999 177654
rect 193397 173906 193463 173909
rect 193673 173906 193739 173909
rect 193397 173904 193739 173906
rect 193397 173848 193402 173904
rect 193458 173848 193678 173904
rect 193734 173848 193739 173904
rect 193397 173846 193739 173848
rect 193397 173843 193463 173846
rect 193673 173843 193739 173846
rect 179505 172546 179571 172549
rect 179689 172546 179755 172549
rect 179505 172544 179755 172546
rect 179505 172488 179510 172544
rect 179566 172488 179694 172544
rect 179750 172488 179755 172544
rect 179505 172486 179755 172488
rect 179505 172483 179571 172486
rect 179689 172483 179755 172486
rect 579889 170098 579955 170101
rect 583520 170098 584960 170188
rect 579889 170096 584960 170098
rect 579889 170040 579894 170096
rect 579950 170040 584960 170096
rect 579889 170038 584960 170040
rect 579889 170035 579955 170038
rect 583520 169948 584960 170038
rect -960 165066 480 165156
rect 3233 165066 3299 165069
rect -960 165064 3299 165066
rect -960 165008 3238 165064
rect 3294 165008 3299 165064
rect -960 165006 3299 165008
rect -960 164916 480 165006
rect 3233 165003 3299 165006
rect 159081 164250 159147 164253
rect 159265 164250 159331 164253
rect 159081 164248 159331 164250
rect 159081 164192 159086 164248
rect 159142 164192 159270 164248
rect 159326 164192 159331 164248
rect 159081 164190 159331 164192
rect 159081 164187 159147 164190
rect 159265 164187 159331 164190
rect 193397 164250 193463 164253
rect 193581 164250 193647 164253
rect 193397 164248 193647 164250
rect 193397 164192 193402 164248
rect 193458 164192 193586 164248
rect 193642 164192 193647 164248
rect 193397 164190 193647 164192
rect 193397 164187 193463 164190
rect 193581 164187 193647 164190
rect 206001 164250 206067 164253
rect 206553 164250 206619 164253
rect 206001 164248 206619 164250
rect 206001 164192 206006 164248
rect 206062 164192 206558 164248
rect 206614 164192 206619 164248
rect 206001 164190 206619 164192
rect 206001 164187 206067 164190
rect 206553 164187 206619 164190
rect 217041 164250 217107 164253
rect 217225 164250 217291 164253
rect 217041 164248 217291 164250
rect 217041 164192 217046 164248
rect 217102 164192 217230 164248
rect 217286 164192 217291 164248
rect 217041 164190 217291 164192
rect 217041 164187 217107 164190
rect 217225 164187 217291 164190
rect 222561 164250 222627 164253
rect 222929 164250 222995 164253
rect 222561 164248 222995 164250
rect 222561 164192 222566 164248
rect 222622 164192 222934 164248
rect 222990 164192 222995 164248
rect 222561 164190 222995 164192
rect 222561 164187 222627 164190
rect 222929 164187 222995 164190
rect 226701 164250 226767 164253
rect 227069 164250 227135 164253
rect 226701 164248 227135 164250
rect 226701 164192 226706 164248
rect 226762 164192 227074 164248
rect 227130 164192 227135 164248
rect 226701 164190 227135 164192
rect 226701 164187 226767 164190
rect 227069 164187 227135 164190
rect 227989 164250 228055 164253
rect 228265 164250 228331 164253
rect 227989 164248 228331 164250
rect 227989 164192 227994 164248
rect 228050 164192 228270 164248
rect 228326 164192 228331 164248
rect 227989 164190 228331 164192
rect 227989 164187 228055 164190
rect 228265 164187 228331 164190
rect 185117 162890 185183 162893
rect 185301 162890 185367 162893
rect 185117 162888 185367 162890
rect 185117 162832 185122 162888
rect 185178 162832 185306 162888
rect 185362 162832 185367 162888
rect 185117 162830 185367 162832
rect 185117 162827 185183 162830
rect 185301 162827 185367 162830
rect 221089 162890 221155 162893
rect 221365 162890 221431 162893
rect 221089 162888 221431 162890
rect 221089 162832 221094 162888
rect 221150 162832 221370 162888
rect 221426 162832 221431 162888
rect 221089 162830 221431 162832
rect 221089 162827 221155 162830
rect 221365 162827 221431 162830
rect 580165 158402 580231 158405
rect 583520 158402 584960 158492
rect 580165 158400 584960 158402
rect 580165 158344 580170 158400
rect 580226 158344 584960 158400
rect 580165 158342 584960 158344
rect 580165 158339 580231 158342
rect 583520 158252 584960 158342
rect 193581 154730 193647 154733
rect 193446 154728 193647 154730
rect 193446 154672 193586 154728
rect 193642 154672 193647 154728
rect 193446 154670 193647 154672
rect 193446 154597 193506 154670
rect 193581 154667 193647 154670
rect 200389 154730 200455 154733
rect 207197 154730 207263 154733
rect 200389 154728 200498 154730
rect 200389 154672 200394 154728
rect 200450 154672 200498 154728
rect 200389 154667 200498 154672
rect 207197 154728 207306 154730
rect 207197 154672 207202 154728
rect 207258 154672 207306 154728
rect 207197 154667 207306 154672
rect 200438 154597 200498 154667
rect 207246 154597 207306 154667
rect 157609 154594 157675 154597
rect 157793 154594 157859 154597
rect 157609 154592 157859 154594
rect 157609 154536 157614 154592
rect 157670 154536 157798 154592
rect 157854 154536 157859 154592
rect 157609 154534 157859 154536
rect 157609 154531 157675 154534
rect 157793 154531 157859 154534
rect 168373 154594 168439 154597
rect 168557 154594 168623 154597
rect 168373 154592 168623 154594
rect 168373 154536 168378 154592
rect 168434 154536 168562 154592
rect 168618 154536 168623 154592
rect 168373 154534 168623 154536
rect 168373 154531 168439 154534
rect 168557 154531 168623 154534
rect 172421 154594 172487 154597
rect 172605 154594 172671 154597
rect 172421 154592 172671 154594
rect 172421 154536 172426 154592
rect 172482 154536 172610 154592
rect 172666 154536 172671 154592
rect 172421 154534 172671 154536
rect 193446 154592 193555 154597
rect 193446 154536 193494 154592
rect 193550 154536 193555 154592
rect 193446 154534 193555 154536
rect 172421 154531 172487 154534
rect 172605 154531 172671 154534
rect 193489 154531 193555 154534
rect 198733 154594 198799 154597
rect 199009 154594 199075 154597
rect 198733 154592 199075 154594
rect 198733 154536 198738 154592
rect 198794 154536 199014 154592
rect 199070 154536 199075 154592
rect 198733 154534 199075 154536
rect 198733 154531 198799 154534
rect 199009 154531 199075 154534
rect 200389 154592 200498 154597
rect 200389 154536 200394 154592
rect 200450 154536 200498 154592
rect 200389 154534 200498 154536
rect 207197 154592 207306 154597
rect 207197 154536 207202 154592
rect 207258 154536 207306 154592
rect 207197 154534 207306 154536
rect 256785 154594 256851 154597
rect 256969 154594 257035 154597
rect 256785 154592 257035 154594
rect 256785 154536 256790 154592
rect 256846 154536 256974 154592
rect 257030 154536 257035 154592
rect 256785 154534 257035 154536
rect 200389 154531 200455 154534
rect 207197 154531 207263 154534
rect 256785 154531 256851 154534
rect 256969 154531 257035 154534
rect 179689 153234 179755 153237
rect 179873 153234 179939 153237
rect 179689 153232 179939 153234
rect 179689 153176 179694 153232
rect 179750 153176 179878 153232
rect 179934 153176 179939 153232
rect 179689 153174 179939 153176
rect 179689 153171 179755 153174
rect 179873 153171 179939 153174
rect -960 150786 480 150876
rect 3693 150786 3759 150789
rect -960 150784 3759 150786
rect -960 150728 3698 150784
rect 3754 150728 3759 150784
rect -960 150726 3759 150728
rect -960 150636 480 150726
rect 3693 150723 3759 150726
rect 583520 146556 584960 146796
rect 157609 145072 157675 145077
rect 158989 145074 159055 145077
rect 157609 145016 157614 145072
rect 157670 145016 157675 145072
rect 157609 145011 157675 145016
rect 158854 145072 159055 145074
rect 158854 145016 158994 145072
rect 159050 145016 159055 145072
rect 158854 145014 159055 145016
rect 157612 144941 157672 145011
rect 157609 144936 157675 144941
rect 157609 144880 157614 144936
rect 157670 144880 157675 144936
rect 157609 144875 157675 144880
rect 158854 144938 158914 145014
rect 158989 145011 159055 145014
rect 198733 145074 198799 145077
rect 217041 145074 217107 145077
rect 198733 145072 198842 145074
rect 198733 145016 198738 145072
rect 198794 145016 198842 145072
rect 198733 145011 198842 145016
rect 158989 144938 159055 144941
rect 158854 144936 159055 144938
rect 158854 144880 158994 144936
rect 159050 144880 159055 144936
rect 158854 144878 159055 144880
rect 158989 144875 159055 144878
rect 194133 144802 194199 144805
rect 198782 144802 198842 145011
rect 216998 145072 217107 145074
rect 216998 145016 217046 145072
rect 217102 145016 217107 145072
rect 216998 145011 217107 145016
rect 216998 144941 217058 145011
rect 216998 144936 217107 144941
rect 216998 144880 217046 144936
rect 217102 144880 217107 144936
rect 216998 144878 217107 144880
rect 217041 144875 217107 144878
rect 256877 144938 256943 144941
rect 257153 144938 257219 144941
rect 256877 144936 257219 144938
rect 256877 144880 256882 144936
rect 256938 144880 257158 144936
rect 257214 144880 257219 144936
rect 256877 144878 257219 144880
rect 256877 144875 256943 144878
rect 257153 144875 257219 144878
rect 194133 144800 198842 144802
rect 194133 144744 194138 144800
rect 194194 144744 198842 144800
rect 194133 144742 198842 144744
rect 194133 144739 194199 144742
rect 163037 143578 163103 143581
rect 163221 143578 163287 143581
rect 163037 143576 163287 143578
rect 163037 143520 163042 143576
rect 163098 143520 163226 143576
rect 163282 143520 163287 143576
rect 163037 143518 163287 143520
rect 163037 143515 163103 143518
rect 163221 143515 163287 143518
rect 225229 143578 225295 143581
rect 225413 143578 225479 143581
rect 225229 143576 225479 143578
rect 225229 143520 225234 143576
rect 225290 143520 225418 143576
rect 225474 143520 225479 143576
rect 225229 143518 225479 143520
rect 225229 143515 225295 143518
rect 225413 143515 225479 143518
rect -960 136370 480 136460
rect 3325 136370 3391 136373
rect -960 136368 3391 136370
rect -960 136312 3330 136368
rect 3386 136312 3391 136368
rect -960 136310 3391 136312
rect -960 136220 480 136310
rect 3325 136307 3391 136310
rect 196249 135418 196315 135421
rect 196206 135416 196315 135418
rect 196206 135360 196254 135416
rect 196310 135360 196315 135416
rect 196206 135355 196315 135360
rect 196206 135285 196266 135355
rect 196157 135280 196266 135285
rect 196157 135224 196162 135280
rect 196218 135224 196266 135280
rect 196157 135222 196266 135224
rect 197629 135282 197695 135285
rect 197813 135282 197879 135285
rect 197629 135280 197879 135282
rect 197629 135224 197634 135280
rect 197690 135224 197818 135280
rect 197874 135224 197879 135280
rect 197629 135222 197879 135224
rect 196157 135219 196223 135222
rect 197629 135219 197695 135222
rect 197813 135219 197879 135222
rect 579889 134874 579955 134877
rect 583520 134874 584960 134964
rect 579889 134872 584960 134874
rect 579889 134816 579894 134872
rect 579950 134816 584960 134872
rect 579889 134814 584960 134816
rect 579889 134811 579955 134814
rect 583520 134724 584960 134814
rect 168373 133922 168439 133925
rect 168557 133922 168623 133925
rect 168373 133920 168623 133922
rect 168373 133864 168378 133920
rect 168434 133864 168562 133920
rect 168618 133864 168623 133920
rect 168373 133862 168623 133864
rect 168373 133859 168439 133862
rect 168557 133859 168623 133862
rect 218237 125626 218303 125629
rect 218421 125626 218487 125629
rect 218237 125624 218487 125626
rect 218237 125568 218242 125624
rect 218298 125568 218426 125624
rect 218482 125568 218487 125624
rect 218237 125566 218487 125568
rect 218237 125563 218303 125566
rect 218421 125563 218487 125566
rect 220997 125626 221063 125629
rect 221181 125626 221247 125629
rect 220997 125624 221247 125626
rect 220997 125568 221002 125624
rect 221058 125568 221186 125624
rect 221242 125568 221247 125624
rect 220997 125566 221247 125568
rect 220997 125563 221063 125566
rect 221181 125563 221247 125566
rect 256877 125626 256943 125629
rect 257153 125626 257219 125629
rect 256877 125624 257219 125626
rect 256877 125568 256882 125624
rect 256938 125568 257158 125624
rect 257214 125568 257219 125624
rect 256877 125566 257219 125568
rect 256877 125563 256943 125566
rect 257153 125563 257219 125566
rect 579889 123178 579955 123181
rect 583520 123178 584960 123268
rect 579889 123176 584960 123178
rect 579889 123120 579894 123176
rect 579950 123120 584960 123176
rect 579889 123118 584960 123120
rect 579889 123115 579955 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 3325 122090 3391 122093
rect -960 122088 3391 122090
rect -960 122032 3330 122088
rect 3386 122032 3391 122088
rect -960 122030 3391 122032
rect -960 121940 480 122030
rect 3325 122027 3391 122030
rect 209865 115970 209931 115973
rect 210141 115970 210207 115973
rect 209865 115968 210207 115970
rect 209865 115912 209870 115968
rect 209926 115912 210146 115968
rect 210202 115912 210207 115968
rect 209865 115910 210207 115912
rect 209865 115907 209931 115910
rect 210141 115907 210207 115910
rect 221089 113250 221155 113253
rect 221273 113250 221339 113253
rect 221089 113248 221339 113250
rect 221089 113192 221094 113248
rect 221150 113192 221278 113248
rect 221334 113192 221339 113248
rect 221089 113190 221339 113192
rect 221089 113187 221155 113190
rect 221273 113187 221339 113190
rect 580165 111482 580231 111485
rect 583520 111482 584960 111572
rect 580165 111480 584960 111482
rect 580165 111424 580170 111480
rect 580226 111424 584960 111480
rect 580165 111422 584960 111424
rect 580165 111419 580231 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3601 107674 3667 107677
rect -960 107672 3667 107674
rect -960 107616 3606 107672
rect 3662 107616 3667 107672
rect -960 107614 3667 107616
rect -960 107524 480 107614
rect 3601 107611 3667 107614
rect 256877 106314 256943 106317
rect 257153 106314 257219 106317
rect 256877 106312 257219 106314
rect 256877 106256 256882 106312
rect 256938 106256 257158 106312
rect 257214 106256 257219 106312
rect 256877 106254 257219 106256
rect 256877 106251 256943 106254
rect 257153 106251 257219 106254
rect 583520 99636 584960 99876
rect 209865 96658 209931 96661
rect 210141 96658 210207 96661
rect 209865 96656 210207 96658
rect 209865 96600 209870 96656
rect 209926 96600 210146 96656
rect 210202 96600 210207 96656
rect 209865 96598 210207 96600
rect 209865 96595 209931 96598
rect 210141 96595 210207 96598
rect -960 93258 480 93348
rect 3601 93258 3667 93261
rect -960 93256 3667 93258
rect -960 93200 3606 93256
rect 3662 93200 3667 93256
rect -960 93198 3667 93200
rect -960 93108 480 93198
rect 3601 93195 3667 93198
rect 579889 87954 579955 87957
rect 583520 87954 584960 88044
rect 579889 87952 584960 87954
rect 579889 87896 579894 87952
rect 579950 87896 584960 87952
rect 579889 87894 584960 87896
rect 579889 87891 579955 87894
rect 583520 87804 584960 87894
rect -960 78978 480 79068
rect 3049 78978 3115 78981
rect -960 78976 3115 78978
rect -960 78920 3054 78976
rect 3110 78920 3115 78976
rect -960 78918 3115 78920
rect -960 78828 480 78918
rect 3049 78915 3115 78918
rect 579889 76258 579955 76261
rect 583520 76258 584960 76348
rect 579889 76256 584960 76258
rect 579889 76200 579894 76256
rect 579950 76200 584960 76256
rect 579889 76198 584960 76200
rect 579889 76195 579955 76198
rect 583520 76108 584960 76198
rect 183921 74762 183987 74765
rect 183694 74760 183987 74762
rect 183694 74704 183926 74760
rect 183982 74704 183987 74760
rect 183694 74702 183987 74704
rect 183694 74626 183754 74702
rect 183921 74699 183987 74702
rect 183829 74626 183895 74629
rect 183694 74624 183895 74626
rect 183694 74568 183834 74624
rect 183890 74568 183895 74624
rect 183694 74566 183895 74568
rect 183829 74563 183895 74566
rect 158713 67690 158779 67693
rect 158989 67690 159055 67693
rect 158713 67688 159055 67690
rect 158713 67632 158718 67688
rect 158774 67632 158994 67688
rect 159050 67632 159055 67688
rect 158713 67630 159055 67632
rect 158713 67627 158779 67630
rect 158989 67627 159055 67630
rect 385033 66196 385099 66197
rect 384982 66132 384988 66196
rect 385052 66194 385099 66196
rect 385052 66192 385144 66194
rect 385094 66136 385144 66192
rect 385052 66134 385144 66136
rect 385052 66132 385099 66134
rect 385033 66131 385099 66132
rect -960 64562 480 64652
rect 3509 64562 3575 64565
rect -960 64560 3575 64562
rect -960 64504 3514 64560
rect 3570 64504 3575 64560
rect -960 64502 3575 64504
rect -960 64412 480 64502
rect 3509 64499 3575 64502
rect 580165 64562 580231 64565
rect 583520 64562 584960 64652
rect 580165 64560 584960 64562
rect 580165 64504 580170 64560
rect 580226 64504 584960 64560
rect 580165 64502 584960 64504
rect 580165 64499 580231 64502
rect 583520 64412 584960 64502
rect 384982 60556 384988 60620
rect 385052 60618 385058 60620
rect 385125 60618 385191 60621
rect 385052 60616 385191 60618
rect 385052 60560 385130 60616
rect 385186 60560 385191 60616
rect 385052 60558 385191 60560
rect 385052 60556 385058 60558
rect 385125 60555 385191 60558
rect 256509 57898 256575 57901
rect 256693 57898 256759 57901
rect 256509 57896 256759 57898
rect 256509 57840 256514 57896
rect 256570 57840 256698 57896
rect 256754 57840 256759 57896
rect 256509 57838 256759 57840
rect 256509 57835 256575 57838
rect 256693 57835 256759 57838
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3049 50146 3115 50149
rect -960 50144 3115 50146
rect -960 50088 3054 50144
rect 3110 50088 3115 50144
rect -960 50086 3115 50088
rect -960 49996 480 50086
rect 3049 50083 3115 50086
rect 579889 41034 579955 41037
rect 583520 41034 584960 41124
rect 579889 41032 584960 41034
rect 579889 40976 579894 41032
rect 579950 40976 584960 41032
rect 579889 40974 584960 40976
rect 579889 40971 579955 40974
rect 583520 40884 584960 40974
rect 256509 38586 256575 38589
rect 256693 38586 256759 38589
rect 256509 38584 256759 38586
rect 256509 38528 256514 38584
rect 256570 38528 256698 38584
rect 256754 38528 256759 38584
rect 256509 38526 256759 38528
rect 256509 38523 256575 38526
rect 256693 38523 256759 38526
rect 207289 37498 207355 37501
rect 207246 37496 207355 37498
rect 207246 37440 207294 37496
rect 207350 37440 207355 37496
rect 207246 37435 207355 37440
rect 207246 37362 207306 37435
rect 207381 37362 207447 37365
rect 207246 37360 207447 37362
rect 207246 37304 207386 37360
rect 207442 37304 207447 37360
rect 207246 37302 207447 37304
rect 207381 37299 207447 37302
rect -960 35866 480 35956
rect 3509 35866 3575 35869
rect -960 35864 3575 35866
rect -960 35808 3514 35864
rect 3570 35808 3575 35864
rect -960 35806 3575 35808
rect -960 35716 480 35806
rect 3509 35803 3575 35806
rect 579889 29338 579955 29341
rect 583520 29338 584960 29428
rect 579889 29336 584960 29338
rect 579889 29280 579894 29336
rect 579950 29280 584960 29336
rect 579889 29278 584960 29280
rect 579889 29275 579955 29278
rect 583520 29188 584960 29278
rect -960 21450 480 21540
rect 3417 21450 3483 21453
rect -960 21448 3483 21450
rect -960 21392 3422 21448
rect 3478 21392 3483 21448
rect -960 21390 3483 21392
rect -960 21300 480 21390
rect 3417 21387 3483 21390
rect 580257 17642 580323 17645
rect 583520 17642 584960 17732
rect 580257 17640 584960 17642
rect 580257 17584 580262 17640
rect 580318 17584 584960 17640
rect 580257 17582 584960 17584
rect 580257 17579 580323 17582
rect 583520 17492 584960 17582
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 583520 5796 584960 6036
rect 20713 3770 20779 3773
rect 162945 3770 163011 3773
rect 20713 3768 163011 3770
rect 20713 3712 20718 3768
rect 20774 3712 162950 3768
rect 163006 3712 163011 3768
rect 20713 3710 163011 3712
rect 20713 3707 20779 3710
rect 162945 3707 163011 3710
rect 299381 3770 299447 3773
rect 357341 3770 357407 3773
rect 299381 3768 357407 3770
rect 299381 3712 299386 3768
rect 299442 3712 357346 3768
rect 357402 3712 357407 3768
rect 299381 3710 357407 3712
rect 299381 3707 299447 3710
rect 357341 3707 357407 3710
rect 382181 3770 382247 3773
rect 564341 3770 564407 3773
rect 382181 3768 564407 3770
rect 382181 3712 382186 3768
rect 382242 3712 564346 3768
rect 564402 3712 564407 3768
rect 382181 3710 564407 3712
rect 382181 3707 382247 3710
rect 564341 3707 564407 3710
rect 19517 3634 19583 3637
rect 162853 3634 162919 3637
rect 19517 3632 162919 3634
rect 19517 3576 19522 3632
rect 19578 3576 162858 3632
rect 162914 3576 162919 3632
rect 19517 3574 162919 3576
rect 19517 3571 19583 3574
rect 162853 3571 162919 3574
rect 302141 3634 302207 3637
rect 364517 3634 364583 3637
rect 302141 3632 364583 3634
rect 302141 3576 302146 3632
rect 302202 3576 364522 3632
rect 364578 3576 364583 3632
rect 302141 3574 364583 3576
rect 302141 3571 302207 3574
rect 364517 3571 364583 3574
rect 386321 3634 386387 3637
rect 571425 3634 571491 3637
rect 386321 3632 571491 3634
rect 386321 3576 386326 3632
rect 386382 3576 571430 3632
rect 571486 3576 571491 3632
rect 386321 3574 571491 3576
rect 386321 3571 386387 3574
rect 571425 3571 571491 3574
rect 11237 3498 11303 3501
rect 158989 3498 159055 3501
rect 11237 3496 159055 3498
rect 11237 3440 11242 3496
rect 11298 3440 158994 3496
rect 159050 3440 159055 3496
rect 11237 3438 159055 3440
rect 11237 3435 11303 3438
rect 158989 3435 159055 3438
rect 303521 3498 303587 3501
rect 368013 3498 368079 3501
rect 303521 3496 368079 3498
rect 303521 3440 303526 3496
rect 303582 3440 368018 3496
rect 368074 3440 368079 3496
rect 303521 3438 368079 3440
rect 303521 3435 303587 3438
rect 368013 3435 368079 3438
rect 387701 3498 387767 3501
rect 575013 3498 575079 3501
rect 387701 3496 575079 3498
rect 387701 3440 387706 3496
rect 387762 3440 575018 3496
rect 575074 3440 575079 3496
rect 387701 3438 575079 3440
rect 387701 3435 387767 3438
rect 575013 3435 575079 3438
rect 5257 3362 5323 3365
rect 156413 3362 156479 3365
rect 5257 3360 156479 3362
rect 5257 3304 5262 3360
rect 5318 3304 156418 3360
rect 156474 3304 156479 3360
rect 5257 3302 156479 3304
rect 5257 3299 5323 3302
rect 156413 3299 156479 3302
rect 306281 3362 306347 3365
rect 375189 3362 375255 3365
rect 306281 3360 375255 3362
rect 306281 3304 306286 3360
rect 306342 3304 375194 3360
rect 375250 3304 375255 3360
rect 306281 3302 375255 3304
rect 306281 3299 306347 3302
rect 375189 3299 375255 3302
rect 389081 3362 389147 3365
rect 578601 3362 578667 3365
rect 389081 3360 578667 3362
rect 389081 3304 389086 3360
rect 389142 3304 578606 3360
rect 578662 3304 578667 3360
rect 389081 3302 578667 3304
rect 389081 3299 389147 3302
rect 578601 3299 578667 3302
<< via3 >>
rect 384988 66192 385052 66196
rect 384988 66136 385038 66192
rect 385038 66136 385052 66192
rect 384988 66132 385052 66136
rect 384988 60556 385052 60620
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 679254 -7976 710862
rect -8576 679018 -8394 679254
rect -8158 679018 -7976 679254
rect -8576 678934 -7976 679018
rect -8576 678698 -8394 678934
rect -8158 678698 -7976 678934
rect -8576 643254 -7976 678698
rect -8576 643018 -8394 643254
rect -8158 643018 -7976 643254
rect -8576 642934 -7976 643018
rect -8576 642698 -8394 642934
rect -8158 642698 -7976 642934
rect -8576 607254 -7976 642698
rect -8576 607018 -8394 607254
rect -8158 607018 -7976 607254
rect -8576 606934 -7976 607018
rect -8576 606698 -8394 606934
rect -8158 606698 -7976 606934
rect -8576 571254 -7976 606698
rect -8576 571018 -8394 571254
rect -8158 571018 -7976 571254
rect -8576 570934 -7976 571018
rect -8576 570698 -8394 570934
rect -8158 570698 -7976 570934
rect -8576 535254 -7976 570698
rect -8576 535018 -8394 535254
rect -8158 535018 -7976 535254
rect -8576 534934 -7976 535018
rect -8576 534698 -8394 534934
rect -8158 534698 -7976 534934
rect -8576 499254 -7976 534698
rect -8576 499018 -8394 499254
rect -8158 499018 -7976 499254
rect -8576 498934 -7976 499018
rect -8576 498698 -8394 498934
rect -8158 498698 -7976 498934
rect -8576 463254 -7976 498698
rect -8576 463018 -8394 463254
rect -8158 463018 -7976 463254
rect -8576 462934 -7976 463018
rect -8576 462698 -8394 462934
rect -8158 462698 -7976 462934
rect -8576 427254 -7976 462698
rect -8576 427018 -8394 427254
rect -8158 427018 -7976 427254
rect -8576 426934 -7976 427018
rect -8576 426698 -8394 426934
rect -8158 426698 -7976 426934
rect -8576 391254 -7976 426698
rect -8576 391018 -8394 391254
rect -8158 391018 -7976 391254
rect -8576 390934 -7976 391018
rect -8576 390698 -8394 390934
rect -8158 390698 -7976 390934
rect -8576 355254 -7976 390698
rect -8576 355018 -8394 355254
rect -8158 355018 -7976 355254
rect -8576 354934 -7976 355018
rect -8576 354698 -8394 354934
rect -8158 354698 -7976 354934
rect -8576 319254 -7976 354698
rect -8576 319018 -8394 319254
rect -8158 319018 -7976 319254
rect -8576 318934 -7976 319018
rect -8576 318698 -8394 318934
rect -8158 318698 -7976 318934
rect -8576 283254 -7976 318698
rect -8576 283018 -8394 283254
rect -8158 283018 -7976 283254
rect -8576 282934 -7976 283018
rect -8576 282698 -8394 282934
rect -8158 282698 -7976 282934
rect -8576 247254 -7976 282698
rect -8576 247018 -8394 247254
rect -8158 247018 -7976 247254
rect -8576 246934 -7976 247018
rect -8576 246698 -8394 246934
rect -8158 246698 -7976 246934
rect -8576 211254 -7976 246698
rect -8576 211018 -8394 211254
rect -8158 211018 -7976 211254
rect -8576 210934 -7976 211018
rect -8576 210698 -8394 210934
rect -8158 210698 -7976 210934
rect -8576 175254 -7976 210698
rect -8576 175018 -8394 175254
rect -8158 175018 -7976 175254
rect -8576 174934 -7976 175018
rect -8576 174698 -8394 174934
rect -8158 174698 -7976 174934
rect -8576 139254 -7976 174698
rect -8576 139018 -8394 139254
rect -8158 139018 -7976 139254
rect -8576 138934 -7976 139018
rect -8576 138698 -8394 138934
rect -8158 138698 -7976 138934
rect -8576 103254 -7976 138698
rect -8576 103018 -8394 103254
rect -8158 103018 -7976 103254
rect -8576 102934 -7976 103018
rect -8576 102698 -8394 102934
rect -8158 102698 -7976 102934
rect -8576 67254 -7976 102698
rect -8576 67018 -8394 67254
rect -8158 67018 -7976 67254
rect -8576 66934 -7976 67018
rect -8576 66698 -8394 66934
rect -8158 66698 -7976 66934
rect -8576 31254 -7976 66698
rect -8576 31018 -8394 31254
rect -8158 31018 -7976 31254
rect -8576 30934 -7976 31018
rect -8576 30698 -8394 30934
rect -8158 30698 -7976 30934
rect -8576 -6926 -7976 30698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 697254 -7036 709922
rect 11604 710478 12204 711440
rect 11604 710242 11786 710478
rect 12022 710242 12204 710478
rect 11604 710158 12204 710242
rect 11604 709922 11786 710158
rect 12022 709922 12204 710158
rect -7636 697018 -7454 697254
rect -7218 697018 -7036 697254
rect -7636 696934 -7036 697018
rect -7636 696698 -7454 696934
rect -7218 696698 -7036 696934
rect -7636 661254 -7036 696698
rect -7636 661018 -7454 661254
rect -7218 661018 -7036 661254
rect -7636 660934 -7036 661018
rect -7636 660698 -7454 660934
rect -7218 660698 -7036 660934
rect -7636 625254 -7036 660698
rect -7636 625018 -7454 625254
rect -7218 625018 -7036 625254
rect -7636 624934 -7036 625018
rect -7636 624698 -7454 624934
rect -7218 624698 -7036 624934
rect -7636 589254 -7036 624698
rect -7636 589018 -7454 589254
rect -7218 589018 -7036 589254
rect -7636 588934 -7036 589018
rect -7636 588698 -7454 588934
rect -7218 588698 -7036 588934
rect -7636 553254 -7036 588698
rect -7636 553018 -7454 553254
rect -7218 553018 -7036 553254
rect -7636 552934 -7036 553018
rect -7636 552698 -7454 552934
rect -7218 552698 -7036 552934
rect -7636 517254 -7036 552698
rect -7636 517018 -7454 517254
rect -7218 517018 -7036 517254
rect -7636 516934 -7036 517018
rect -7636 516698 -7454 516934
rect -7218 516698 -7036 516934
rect -7636 481254 -7036 516698
rect -7636 481018 -7454 481254
rect -7218 481018 -7036 481254
rect -7636 480934 -7036 481018
rect -7636 480698 -7454 480934
rect -7218 480698 -7036 480934
rect -7636 445254 -7036 480698
rect -7636 445018 -7454 445254
rect -7218 445018 -7036 445254
rect -7636 444934 -7036 445018
rect -7636 444698 -7454 444934
rect -7218 444698 -7036 444934
rect -7636 409254 -7036 444698
rect -7636 409018 -7454 409254
rect -7218 409018 -7036 409254
rect -7636 408934 -7036 409018
rect -7636 408698 -7454 408934
rect -7218 408698 -7036 408934
rect -7636 373254 -7036 408698
rect -7636 373018 -7454 373254
rect -7218 373018 -7036 373254
rect -7636 372934 -7036 373018
rect -7636 372698 -7454 372934
rect -7218 372698 -7036 372934
rect -7636 337254 -7036 372698
rect -7636 337018 -7454 337254
rect -7218 337018 -7036 337254
rect -7636 336934 -7036 337018
rect -7636 336698 -7454 336934
rect -7218 336698 -7036 336934
rect -7636 301254 -7036 336698
rect -7636 301018 -7454 301254
rect -7218 301018 -7036 301254
rect -7636 300934 -7036 301018
rect -7636 300698 -7454 300934
rect -7218 300698 -7036 300934
rect -7636 265254 -7036 300698
rect -7636 265018 -7454 265254
rect -7218 265018 -7036 265254
rect -7636 264934 -7036 265018
rect -7636 264698 -7454 264934
rect -7218 264698 -7036 264934
rect -7636 229254 -7036 264698
rect -7636 229018 -7454 229254
rect -7218 229018 -7036 229254
rect -7636 228934 -7036 229018
rect -7636 228698 -7454 228934
rect -7218 228698 -7036 228934
rect -7636 193254 -7036 228698
rect -7636 193018 -7454 193254
rect -7218 193018 -7036 193254
rect -7636 192934 -7036 193018
rect -7636 192698 -7454 192934
rect -7218 192698 -7036 192934
rect -7636 157254 -7036 192698
rect -7636 157018 -7454 157254
rect -7218 157018 -7036 157254
rect -7636 156934 -7036 157018
rect -7636 156698 -7454 156934
rect -7218 156698 -7036 156934
rect -7636 121254 -7036 156698
rect -7636 121018 -7454 121254
rect -7218 121018 -7036 121254
rect -7636 120934 -7036 121018
rect -7636 120698 -7454 120934
rect -7218 120698 -7036 120934
rect -7636 85254 -7036 120698
rect -7636 85018 -7454 85254
rect -7218 85018 -7036 85254
rect -7636 84934 -7036 85018
rect -7636 84698 -7454 84934
rect -7218 84698 -7036 84934
rect -7636 49254 -7036 84698
rect -7636 49018 -7454 49254
rect -7218 49018 -7036 49254
rect -7636 48934 -7036 49018
rect -7636 48698 -7454 48934
rect -7218 48698 -7036 48934
rect -7636 13254 -7036 48698
rect -7636 13018 -7454 13254
rect -7218 13018 -7036 13254
rect -7636 12934 -7036 13018
rect -7636 12698 -7454 12934
rect -7218 12698 -7036 12934
rect -7636 -5986 -7036 12698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 675654 -6096 708982
rect -6696 675418 -6514 675654
rect -6278 675418 -6096 675654
rect -6696 675334 -6096 675418
rect -6696 675098 -6514 675334
rect -6278 675098 -6096 675334
rect -6696 639654 -6096 675098
rect -6696 639418 -6514 639654
rect -6278 639418 -6096 639654
rect -6696 639334 -6096 639418
rect -6696 639098 -6514 639334
rect -6278 639098 -6096 639334
rect -6696 603654 -6096 639098
rect -6696 603418 -6514 603654
rect -6278 603418 -6096 603654
rect -6696 603334 -6096 603418
rect -6696 603098 -6514 603334
rect -6278 603098 -6096 603334
rect -6696 567654 -6096 603098
rect -6696 567418 -6514 567654
rect -6278 567418 -6096 567654
rect -6696 567334 -6096 567418
rect -6696 567098 -6514 567334
rect -6278 567098 -6096 567334
rect -6696 531654 -6096 567098
rect -6696 531418 -6514 531654
rect -6278 531418 -6096 531654
rect -6696 531334 -6096 531418
rect -6696 531098 -6514 531334
rect -6278 531098 -6096 531334
rect -6696 495654 -6096 531098
rect -6696 495418 -6514 495654
rect -6278 495418 -6096 495654
rect -6696 495334 -6096 495418
rect -6696 495098 -6514 495334
rect -6278 495098 -6096 495334
rect -6696 459654 -6096 495098
rect -6696 459418 -6514 459654
rect -6278 459418 -6096 459654
rect -6696 459334 -6096 459418
rect -6696 459098 -6514 459334
rect -6278 459098 -6096 459334
rect -6696 423654 -6096 459098
rect -6696 423418 -6514 423654
rect -6278 423418 -6096 423654
rect -6696 423334 -6096 423418
rect -6696 423098 -6514 423334
rect -6278 423098 -6096 423334
rect -6696 387654 -6096 423098
rect -6696 387418 -6514 387654
rect -6278 387418 -6096 387654
rect -6696 387334 -6096 387418
rect -6696 387098 -6514 387334
rect -6278 387098 -6096 387334
rect -6696 351654 -6096 387098
rect -6696 351418 -6514 351654
rect -6278 351418 -6096 351654
rect -6696 351334 -6096 351418
rect -6696 351098 -6514 351334
rect -6278 351098 -6096 351334
rect -6696 315654 -6096 351098
rect -6696 315418 -6514 315654
rect -6278 315418 -6096 315654
rect -6696 315334 -6096 315418
rect -6696 315098 -6514 315334
rect -6278 315098 -6096 315334
rect -6696 279654 -6096 315098
rect -6696 279418 -6514 279654
rect -6278 279418 -6096 279654
rect -6696 279334 -6096 279418
rect -6696 279098 -6514 279334
rect -6278 279098 -6096 279334
rect -6696 243654 -6096 279098
rect -6696 243418 -6514 243654
rect -6278 243418 -6096 243654
rect -6696 243334 -6096 243418
rect -6696 243098 -6514 243334
rect -6278 243098 -6096 243334
rect -6696 207654 -6096 243098
rect -6696 207418 -6514 207654
rect -6278 207418 -6096 207654
rect -6696 207334 -6096 207418
rect -6696 207098 -6514 207334
rect -6278 207098 -6096 207334
rect -6696 171654 -6096 207098
rect -6696 171418 -6514 171654
rect -6278 171418 -6096 171654
rect -6696 171334 -6096 171418
rect -6696 171098 -6514 171334
rect -6278 171098 -6096 171334
rect -6696 135654 -6096 171098
rect -6696 135418 -6514 135654
rect -6278 135418 -6096 135654
rect -6696 135334 -6096 135418
rect -6696 135098 -6514 135334
rect -6278 135098 -6096 135334
rect -6696 99654 -6096 135098
rect -6696 99418 -6514 99654
rect -6278 99418 -6096 99654
rect -6696 99334 -6096 99418
rect -6696 99098 -6514 99334
rect -6278 99098 -6096 99334
rect -6696 63654 -6096 99098
rect -6696 63418 -6514 63654
rect -6278 63418 -6096 63654
rect -6696 63334 -6096 63418
rect -6696 63098 -6514 63334
rect -6278 63098 -6096 63334
rect -6696 27654 -6096 63098
rect -6696 27418 -6514 27654
rect -6278 27418 -6096 27654
rect -6696 27334 -6096 27418
rect -6696 27098 -6514 27334
rect -6278 27098 -6096 27334
rect -6696 -5046 -6096 27098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 693654 -5156 708042
rect 8004 708598 8604 709560
rect 8004 708362 8186 708598
rect 8422 708362 8604 708598
rect 8004 708278 8604 708362
rect 8004 708042 8186 708278
rect 8422 708042 8604 708278
rect -5756 693418 -5574 693654
rect -5338 693418 -5156 693654
rect -5756 693334 -5156 693418
rect -5756 693098 -5574 693334
rect -5338 693098 -5156 693334
rect -5756 657654 -5156 693098
rect -5756 657418 -5574 657654
rect -5338 657418 -5156 657654
rect -5756 657334 -5156 657418
rect -5756 657098 -5574 657334
rect -5338 657098 -5156 657334
rect -5756 621654 -5156 657098
rect -5756 621418 -5574 621654
rect -5338 621418 -5156 621654
rect -5756 621334 -5156 621418
rect -5756 621098 -5574 621334
rect -5338 621098 -5156 621334
rect -5756 585654 -5156 621098
rect -5756 585418 -5574 585654
rect -5338 585418 -5156 585654
rect -5756 585334 -5156 585418
rect -5756 585098 -5574 585334
rect -5338 585098 -5156 585334
rect -5756 549654 -5156 585098
rect -5756 549418 -5574 549654
rect -5338 549418 -5156 549654
rect -5756 549334 -5156 549418
rect -5756 549098 -5574 549334
rect -5338 549098 -5156 549334
rect -5756 513654 -5156 549098
rect -5756 513418 -5574 513654
rect -5338 513418 -5156 513654
rect -5756 513334 -5156 513418
rect -5756 513098 -5574 513334
rect -5338 513098 -5156 513334
rect -5756 477654 -5156 513098
rect -5756 477418 -5574 477654
rect -5338 477418 -5156 477654
rect -5756 477334 -5156 477418
rect -5756 477098 -5574 477334
rect -5338 477098 -5156 477334
rect -5756 441654 -5156 477098
rect -5756 441418 -5574 441654
rect -5338 441418 -5156 441654
rect -5756 441334 -5156 441418
rect -5756 441098 -5574 441334
rect -5338 441098 -5156 441334
rect -5756 405654 -5156 441098
rect -5756 405418 -5574 405654
rect -5338 405418 -5156 405654
rect -5756 405334 -5156 405418
rect -5756 405098 -5574 405334
rect -5338 405098 -5156 405334
rect -5756 369654 -5156 405098
rect -5756 369418 -5574 369654
rect -5338 369418 -5156 369654
rect -5756 369334 -5156 369418
rect -5756 369098 -5574 369334
rect -5338 369098 -5156 369334
rect -5756 333654 -5156 369098
rect -5756 333418 -5574 333654
rect -5338 333418 -5156 333654
rect -5756 333334 -5156 333418
rect -5756 333098 -5574 333334
rect -5338 333098 -5156 333334
rect -5756 297654 -5156 333098
rect -5756 297418 -5574 297654
rect -5338 297418 -5156 297654
rect -5756 297334 -5156 297418
rect -5756 297098 -5574 297334
rect -5338 297098 -5156 297334
rect -5756 261654 -5156 297098
rect -5756 261418 -5574 261654
rect -5338 261418 -5156 261654
rect -5756 261334 -5156 261418
rect -5756 261098 -5574 261334
rect -5338 261098 -5156 261334
rect -5756 225654 -5156 261098
rect -5756 225418 -5574 225654
rect -5338 225418 -5156 225654
rect -5756 225334 -5156 225418
rect -5756 225098 -5574 225334
rect -5338 225098 -5156 225334
rect -5756 189654 -5156 225098
rect -5756 189418 -5574 189654
rect -5338 189418 -5156 189654
rect -5756 189334 -5156 189418
rect -5756 189098 -5574 189334
rect -5338 189098 -5156 189334
rect -5756 153654 -5156 189098
rect -5756 153418 -5574 153654
rect -5338 153418 -5156 153654
rect -5756 153334 -5156 153418
rect -5756 153098 -5574 153334
rect -5338 153098 -5156 153334
rect -5756 117654 -5156 153098
rect -5756 117418 -5574 117654
rect -5338 117418 -5156 117654
rect -5756 117334 -5156 117418
rect -5756 117098 -5574 117334
rect -5338 117098 -5156 117334
rect -5756 81654 -5156 117098
rect -5756 81418 -5574 81654
rect -5338 81418 -5156 81654
rect -5756 81334 -5156 81418
rect -5756 81098 -5574 81334
rect -5338 81098 -5156 81334
rect -5756 45654 -5156 81098
rect -5756 45418 -5574 45654
rect -5338 45418 -5156 45654
rect -5756 45334 -5156 45418
rect -5756 45098 -5574 45334
rect -5338 45098 -5156 45334
rect -5756 9654 -5156 45098
rect -5756 9418 -5574 9654
rect -5338 9418 -5156 9654
rect -5756 9334 -5156 9418
rect -5756 9098 -5574 9334
rect -5338 9098 -5156 9334
rect -5756 -4106 -5156 9098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 672054 -4216 707102
rect -4816 671818 -4634 672054
rect -4398 671818 -4216 672054
rect -4816 671734 -4216 671818
rect -4816 671498 -4634 671734
rect -4398 671498 -4216 671734
rect -4816 636054 -4216 671498
rect -4816 635818 -4634 636054
rect -4398 635818 -4216 636054
rect -4816 635734 -4216 635818
rect -4816 635498 -4634 635734
rect -4398 635498 -4216 635734
rect -4816 600054 -4216 635498
rect -4816 599818 -4634 600054
rect -4398 599818 -4216 600054
rect -4816 599734 -4216 599818
rect -4816 599498 -4634 599734
rect -4398 599498 -4216 599734
rect -4816 564054 -4216 599498
rect -4816 563818 -4634 564054
rect -4398 563818 -4216 564054
rect -4816 563734 -4216 563818
rect -4816 563498 -4634 563734
rect -4398 563498 -4216 563734
rect -4816 528054 -4216 563498
rect -4816 527818 -4634 528054
rect -4398 527818 -4216 528054
rect -4816 527734 -4216 527818
rect -4816 527498 -4634 527734
rect -4398 527498 -4216 527734
rect -4816 492054 -4216 527498
rect -4816 491818 -4634 492054
rect -4398 491818 -4216 492054
rect -4816 491734 -4216 491818
rect -4816 491498 -4634 491734
rect -4398 491498 -4216 491734
rect -4816 456054 -4216 491498
rect -4816 455818 -4634 456054
rect -4398 455818 -4216 456054
rect -4816 455734 -4216 455818
rect -4816 455498 -4634 455734
rect -4398 455498 -4216 455734
rect -4816 420054 -4216 455498
rect -4816 419818 -4634 420054
rect -4398 419818 -4216 420054
rect -4816 419734 -4216 419818
rect -4816 419498 -4634 419734
rect -4398 419498 -4216 419734
rect -4816 384054 -4216 419498
rect -4816 383818 -4634 384054
rect -4398 383818 -4216 384054
rect -4816 383734 -4216 383818
rect -4816 383498 -4634 383734
rect -4398 383498 -4216 383734
rect -4816 348054 -4216 383498
rect -4816 347818 -4634 348054
rect -4398 347818 -4216 348054
rect -4816 347734 -4216 347818
rect -4816 347498 -4634 347734
rect -4398 347498 -4216 347734
rect -4816 312054 -4216 347498
rect -4816 311818 -4634 312054
rect -4398 311818 -4216 312054
rect -4816 311734 -4216 311818
rect -4816 311498 -4634 311734
rect -4398 311498 -4216 311734
rect -4816 276054 -4216 311498
rect -4816 275818 -4634 276054
rect -4398 275818 -4216 276054
rect -4816 275734 -4216 275818
rect -4816 275498 -4634 275734
rect -4398 275498 -4216 275734
rect -4816 240054 -4216 275498
rect -4816 239818 -4634 240054
rect -4398 239818 -4216 240054
rect -4816 239734 -4216 239818
rect -4816 239498 -4634 239734
rect -4398 239498 -4216 239734
rect -4816 204054 -4216 239498
rect -4816 203818 -4634 204054
rect -4398 203818 -4216 204054
rect -4816 203734 -4216 203818
rect -4816 203498 -4634 203734
rect -4398 203498 -4216 203734
rect -4816 168054 -4216 203498
rect -4816 167818 -4634 168054
rect -4398 167818 -4216 168054
rect -4816 167734 -4216 167818
rect -4816 167498 -4634 167734
rect -4398 167498 -4216 167734
rect -4816 132054 -4216 167498
rect -4816 131818 -4634 132054
rect -4398 131818 -4216 132054
rect -4816 131734 -4216 131818
rect -4816 131498 -4634 131734
rect -4398 131498 -4216 131734
rect -4816 96054 -4216 131498
rect -4816 95818 -4634 96054
rect -4398 95818 -4216 96054
rect -4816 95734 -4216 95818
rect -4816 95498 -4634 95734
rect -4398 95498 -4216 95734
rect -4816 60054 -4216 95498
rect -4816 59818 -4634 60054
rect -4398 59818 -4216 60054
rect -4816 59734 -4216 59818
rect -4816 59498 -4634 59734
rect -4398 59498 -4216 59734
rect -4816 24054 -4216 59498
rect -4816 23818 -4634 24054
rect -4398 23818 -4216 24054
rect -4816 23734 -4216 23818
rect -4816 23498 -4634 23734
rect -4398 23498 -4216 23734
rect -4816 -3166 -4216 23498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 690054 -3276 706162
rect 4404 706718 5004 707680
rect 4404 706482 4586 706718
rect 4822 706482 5004 706718
rect 4404 706398 5004 706482
rect 4404 706162 4586 706398
rect 4822 706162 5004 706398
rect -3876 689818 -3694 690054
rect -3458 689818 -3276 690054
rect -3876 689734 -3276 689818
rect -3876 689498 -3694 689734
rect -3458 689498 -3276 689734
rect -3876 654054 -3276 689498
rect -3876 653818 -3694 654054
rect -3458 653818 -3276 654054
rect -3876 653734 -3276 653818
rect -3876 653498 -3694 653734
rect -3458 653498 -3276 653734
rect -3876 618054 -3276 653498
rect -3876 617818 -3694 618054
rect -3458 617818 -3276 618054
rect -3876 617734 -3276 617818
rect -3876 617498 -3694 617734
rect -3458 617498 -3276 617734
rect -3876 582054 -3276 617498
rect -3876 581818 -3694 582054
rect -3458 581818 -3276 582054
rect -3876 581734 -3276 581818
rect -3876 581498 -3694 581734
rect -3458 581498 -3276 581734
rect -3876 546054 -3276 581498
rect -3876 545818 -3694 546054
rect -3458 545818 -3276 546054
rect -3876 545734 -3276 545818
rect -3876 545498 -3694 545734
rect -3458 545498 -3276 545734
rect -3876 510054 -3276 545498
rect -3876 509818 -3694 510054
rect -3458 509818 -3276 510054
rect -3876 509734 -3276 509818
rect -3876 509498 -3694 509734
rect -3458 509498 -3276 509734
rect -3876 474054 -3276 509498
rect -3876 473818 -3694 474054
rect -3458 473818 -3276 474054
rect -3876 473734 -3276 473818
rect -3876 473498 -3694 473734
rect -3458 473498 -3276 473734
rect -3876 438054 -3276 473498
rect -3876 437818 -3694 438054
rect -3458 437818 -3276 438054
rect -3876 437734 -3276 437818
rect -3876 437498 -3694 437734
rect -3458 437498 -3276 437734
rect -3876 402054 -3276 437498
rect -3876 401818 -3694 402054
rect -3458 401818 -3276 402054
rect -3876 401734 -3276 401818
rect -3876 401498 -3694 401734
rect -3458 401498 -3276 401734
rect -3876 366054 -3276 401498
rect -3876 365818 -3694 366054
rect -3458 365818 -3276 366054
rect -3876 365734 -3276 365818
rect -3876 365498 -3694 365734
rect -3458 365498 -3276 365734
rect -3876 330054 -3276 365498
rect -3876 329818 -3694 330054
rect -3458 329818 -3276 330054
rect -3876 329734 -3276 329818
rect -3876 329498 -3694 329734
rect -3458 329498 -3276 329734
rect -3876 294054 -3276 329498
rect -3876 293818 -3694 294054
rect -3458 293818 -3276 294054
rect -3876 293734 -3276 293818
rect -3876 293498 -3694 293734
rect -3458 293498 -3276 293734
rect -3876 258054 -3276 293498
rect -3876 257818 -3694 258054
rect -3458 257818 -3276 258054
rect -3876 257734 -3276 257818
rect -3876 257498 -3694 257734
rect -3458 257498 -3276 257734
rect -3876 222054 -3276 257498
rect -3876 221818 -3694 222054
rect -3458 221818 -3276 222054
rect -3876 221734 -3276 221818
rect -3876 221498 -3694 221734
rect -3458 221498 -3276 221734
rect -3876 186054 -3276 221498
rect -3876 185818 -3694 186054
rect -3458 185818 -3276 186054
rect -3876 185734 -3276 185818
rect -3876 185498 -3694 185734
rect -3458 185498 -3276 185734
rect -3876 150054 -3276 185498
rect -3876 149818 -3694 150054
rect -3458 149818 -3276 150054
rect -3876 149734 -3276 149818
rect -3876 149498 -3694 149734
rect -3458 149498 -3276 149734
rect -3876 114054 -3276 149498
rect -3876 113818 -3694 114054
rect -3458 113818 -3276 114054
rect -3876 113734 -3276 113818
rect -3876 113498 -3694 113734
rect -3458 113498 -3276 113734
rect -3876 78054 -3276 113498
rect -3876 77818 -3694 78054
rect -3458 77818 -3276 78054
rect -3876 77734 -3276 77818
rect -3876 77498 -3694 77734
rect -3458 77498 -3276 77734
rect -3876 42054 -3276 77498
rect -3876 41818 -3694 42054
rect -3458 41818 -3276 42054
rect -3876 41734 -3276 41818
rect -3876 41498 -3694 41734
rect -3458 41498 -3276 41734
rect -3876 6054 -3276 41498
rect -3876 5818 -3694 6054
rect -3458 5818 -3276 6054
rect -3876 5734 -3276 5818
rect -3876 5498 -3694 5734
rect -3458 5498 -3276 5734
rect -3876 -2226 -3276 5498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 4404 690054 5004 706162
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 4404 -2226 5004 5498
rect 4404 -2462 4586 -2226
rect 4822 -2462 5004 -2226
rect 4404 -2546 5004 -2462
rect 4404 -2782 4586 -2546
rect 4822 -2782 5004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 4404 -3744 5004 -2782
rect 8004 693654 8604 708042
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 8004 -4106 8604 9098
rect 8004 -4342 8186 -4106
rect 8422 -4342 8604 -4106
rect 8004 -4426 8604 -4342
rect 8004 -4662 8186 -4426
rect 8422 -4662 8604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 8004 -5624 8604 -4662
rect 11604 697254 12204 709922
rect 29604 711418 30204 711440
rect 29604 711182 29786 711418
rect 30022 711182 30204 711418
rect 29604 711098 30204 711182
rect 29604 710862 29786 711098
rect 30022 710862 30204 711098
rect 26004 709538 26604 709560
rect 26004 709302 26186 709538
rect 26422 709302 26604 709538
rect 26004 709218 26604 709302
rect 26004 708982 26186 709218
rect 26422 708982 26604 709218
rect 22404 707658 23004 707680
rect 22404 707422 22586 707658
rect 22822 707422 23004 707658
rect 22404 707338 23004 707422
rect 22404 707102 22586 707338
rect 22822 707102 23004 707338
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 11604 -5986 12204 12698
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 22404 672054 23004 707102
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3166 23004 23498
rect 22404 -3402 22586 -3166
rect 22822 -3402 23004 -3166
rect 22404 -3486 23004 -3402
rect 22404 -3722 22586 -3486
rect 22822 -3722 23004 -3486
rect 22404 -3744 23004 -3722
rect 26004 675654 26604 708982
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -5046 26604 27098
rect 26004 -5282 26186 -5046
rect 26422 -5282 26604 -5046
rect 26004 -5366 26604 -5282
rect 26004 -5602 26186 -5366
rect 26422 -5602 26604 -5366
rect 26004 -5624 26604 -5602
rect 29604 679254 30204 710862
rect 47604 710478 48204 711440
rect 47604 710242 47786 710478
rect 48022 710242 48204 710478
rect 47604 710158 48204 710242
rect 47604 709922 47786 710158
rect 48022 709922 48204 710158
rect 44004 708598 44604 709560
rect 44004 708362 44186 708598
rect 44422 708362 44604 708598
rect 44004 708278 44604 708362
rect 44004 708042 44186 708278
rect 44422 708042 44604 708278
rect 40404 706718 41004 707680
rect 40404 706482 40586 706718
rect 40822 706482 41004 706718
rect 40404 706398 41004 706482
rect 40404 706162 40586 706398
rect 40822 706162 41004 706398
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6222 11786 -5986
rect 12022 -6222 12204 -5986
rect 11604 -6306 12204 -6222
rect 11604 -6542 11786 -6306
rect 12022 -6542 12204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 11604 -7504 12204 -6542
rect 29604 -6926 30204 30698
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 40404 690054 41004 706162
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2226 41004 5498
rect 40404 -2462 40586 -2226
rect 40822 -2462 41004 -2226
rect 40404 -2546 41004 -2462
rect 40404 -2782 40586 -2546
rect 40822 -2782 41004 -2546
rect 40404 -3744 41004 -2782
rect 44004 693654 44604 708042
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4106 44604 9098
rect 44004 -4342 44186 -4106
rect 44422 -4342 44604 -4106
rect 44004 -4426 44604 -4342
rect 44004 -4662 44186 -4426
rect 44422 -4662 44604 -4426
rect 44004 -5624 44604 -4662
rect 47604 697254 48204 709922
rect 65604 711418 66204 711440
rect 65604 711182 65786 711418
rect 66022 711182 66204 711418
rect 65604 711098 66204 711182
rect 65604 710862 65786 711098
rect 66022 710862 66204 711098
rect 62004 709538 62604 709560
rect 62004 709302 62186 709538
rect 62422 709302 62604 709538
rect 62004 709218 62604 709302
rect 62004 708982 62186 709218
rect 62422 708982 62604 709218
rect 58404 707658 59004 707680
rect 58404 707422 58586 707658
rect 58822 707422 59004 707658
rect 58404 707338 59004 707422
rect 58404 707102 58586 707338
rect 58822 707102 59004 707338
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7162 29786 -6926
rect 30022 -7162 30204 -6926
rect 29604 -7246 30204 -7162
rect 29604 -7482 29786 -7246
rect 30022 -7482 30204 -7246
rect 29604 -7504 30204 -7482
rect 47604 -5986 48204 12698
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 58404 672054 59004 707102
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3166 59004 23498
rect 58404 -3402 58586 -3166
rect 58822 -3402 59004 -3166
rect 58404 -3486 59004 -3402
rect 58404 -3722 58586 -3486
rect 58822 -3722 59004 -3486
rect 58404 -3744 59004 -3722
rect 62004 675654 62604 708982
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -5046 62604 27098
rect 62004 -5282 62186 -5046
rect 62422 -5282 62604 -5046
rect 62004 -5366 62604 -5282
rect 62004 -5602 62186 -5366
rect 62422 -5602 62604 -5366
rect 62004 -5624 62604 -5602
rect 65604 679254 66204 710862
rect 83604 710478 84204 711440
rect 83604 710242 83786 710478
rect 84022 710242 84204 710478
rect 83604 710158 84204 710242
rect 83604 709922 83786 710158
rect 84022 709922 84204 710158
rect 80004 708598 80604 709560
rect 80004 708362 80186 708598
rect 80422 708362 80604 708598
rect 80004 708278 80604 708362
rect 80004 708042 80186 708278
rect 80422 708042 80604 708278
rect 76404 706718 77004 707680
rect 76404 706482 76586 706718
rect 76822 706482 77004 706718
rect 76404 706398 77004 706482
rect 76404 706162 76586 706398
rect 76822 706162 77004 706398
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6222 47786 -5986
rect 48022 -6222 48204 -5986
rect 47604 -6306 48204 -6222
rect 47604 -6542 47786 -6306
rect 48022 -6542 48204 -6306
rect 47604 -7504 48204 -6542
rect 65604 -6926 66204 30698
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 76404 690054 77004 706162
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2226 77004 5498
rect 76404 -2462 76586 -2226
rect 76822 -2462 77004 -2226
rect 76404 -2546 77004 -2462
rect 76404 -2782 76586 -2546
rect 76822 -2782 77004 -2546
rect 76404 -3744 77004 -2782
rect 80004 693654 80604 708042
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4106 80604 9098
rect 80004 -4342 80186 -4106
rect 80422 -4342 80604 -4106
rect 80004 -4426 80604 -4342
rect 80004 -4662 80186 -4426
rect 80422 -4662 80604 -4426
rect 80004 -5624 80604 -4662
rect 83604 697254 84204 709922
rect 101604 711418 102204 711440
rect 101604 711182 101786 711418
rect 102022 711182 102204 711418
rect 101604 711098 102204 711182
rect 101604 710862 101786 711098
rect 102022 710862 102204 711098
rect 98004 709538 98604 709560
rect 98004 709302 98186 709538
rect 98422 709302 98604 709538
rect 98004 709218 98604 709302
rect 98004 708982 98186 709218
rect 98422 708982 98604 709218
rect 94404 707658 95004 707680
rect 94404 707422 94586 707658
rect 94822 707422 95004 707658
rect 94404 707338 95004 707422
rect 94404 707102 94586 707338
rect 94822 707102 95004 707338
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 373254 84204 408698
rect 83604 373018 83786 373254
rect 84022 373018 84204 373254
rect 83604 372934 84204 373018
rect 83604 372698 83786 372934
rect 84022 372698 84204 372934
rect 83604 337254 84204 372698
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7162 65786 -6926
rect 66022 -7162 66204 -6926
rect 65604 -7246 66204 -7162
rect 65604 -7482 65786 -7246
rect 66022 -7482 66204 -7246
rect 65604 -7504 66204 -7482
rect 83604 -5986 84204 12698
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 94404 672054 95004 707102
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3166 95004 23498
rect 94404 -3402 94586 -3166
rect 94822 -3402 95004 -3166
rect 94404 -3486 95004 -3402
rect 94404 -3722 94586 -3486
rect 94822 -3722 95004 -3486
rect 94404 -3744 95004 -3722
rect 98004 675654 98604 708982
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 531654 98604 567098
rect 98004 531418 98186 531654
rect 98422 531418 98604 531654
rect 98004 531334 98604 531418
rect 98004 531098 98186 531334
rect 98422 531098 98604 531334
rect 98004 495654 98604 531098
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 387654 98604 423098
rect 98004 387418 98186 387654
rect 98422 387418 98604 387654
rect 98004 387334 98604 387418
rect 98004 387098 98186 387334
rect 98422 387098 98604 387334
rect 98004 351654 98604 387098
rect 98004 351418 98186 351654
rect 98422 351418 98604 351654
rect 98004 351334 98604 351418
rect 98004 351098 98186 351334
rect 98422 351098 98604 351334
rect 98004 315654 98604 351098
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -5046 98604 27098
rect 98004 -5282 98186 -5046
rect 98422 -5282 98604 -5046
rect 98004 -5366 98604 -5282
rect 98004 -5602 98186 -5366
rect 98422 -5602 98604 -5366
rect 98004 -5624 98604 -5602
rect 101604 679254 102204 710862
rect 119604 710478 120204 711440
rect 119604 710242 119786 710478
rect 120022 710242 120204 710478
rect 119604 710158 120204 710242
rect 119604 709922 119786 710158
rect 120022 709922 120204 710158
rect 116004 708598 116604 709560
rect 116004 708362 116186 708598
rect 116422 708362 116604 708598
rect 116004 708278 116604 708362
rect 116004 708042 116186 708278
rect 116422 708042 116604 708278
rect 112404 706718 113004 707680
rect 112404 706482 112586 706718
rect 112822 706482 113004 706718
rect 112404 706398 113004 706482
rect 112404 706162 112586 706398
rect 112822 706162 113004 706398
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 535254 102204 570698
rect 101604 535018 101786 535254
rect 102022 535018 102204 535254
rect 101604 534934 102204 535018
rect 101604 534698 101786 534934
rect 102022 534698 102204 534934
rect 101604 499254 102204 534698
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 391254 102204 426698
rect 101604 391018 101786 391254
rect 102022 391018 102204 391254
rect 101604 390934 102204 391018
rect 101604 390698 101786 390934
rect 102022 390698 102204 390934
rect 101604 355254 102204 390698
rect 101604 355018 101786 355254
rect 102022 355018 102204 355254
rect 101604 354934 102204 355018
rect 101604 354698 101786 354934
rect 102022 354698 102204 354934
rect 101604 319254 102204 354698
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6222 83786 -5986
rect 84022 -6222 84204 -5986
rect 83604 -6306 84204 -6222
rect 83604 -6542 83786 -6306
rect 84022 -6542 84204 -6306
rect 83604 -7504 84204 -6542
rect 101604 -6926 102204 30698
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 112404 690054 113004 706162
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2226 113004 5498
rect 112404 -2462 112586 -2226
rect 112822 -2462 113004 -2226
rect 112404 -2546 113004 -2462
rect 112404 -2782 112586 -2546
rect 112822 -2782 113004 -2546
rect 112404 -3744 113004 -2782
rect 116004 693654 116604 708042
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 369654 116604 405098
rect 116004 369418 116186 369654
rect 116422 369418 116604 369654
rect 116004 369334 116604 369418
rect 116004 369098 116186 369334
rect 116422 369098 116604 369334
rect 116004 333654 116604 369098
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4106 116604 9098
rect 116004 -4342 116186 -4106
rect 116422 -4342 116604 -4106
rect 116004 -4426 116604 -4342
rect 116004 -4662 116186 -4426
rect 116422 -4662 116604 -4426
rect 116004 -5624 116604 -4662
rect 119604 697254 120204 709922
rect 137604 711418 138204 711440
rect 137604 711182 137786 711418
rect 138022 711182 138204 711418
rect 137604 711098 138204 711182
rect 137604 710862 137786 711098
rect 138022 710862 138204 711098
rect 134004 709538 134604 709560
rect 134004 709302 134186 709538
rect 134422 709302 134604 709538
rect 134004 709218 134604 709302
rect 134004 708982 134186 709218
rect 134422 708982 134604 709218
rect 130404 707658 131004 707680
rect 130404 707422 130586 707658
rect 130822 707422 131004 707658
rect 130404 707338 131004 707422
rect 130404 707102 130586 707338
rect 130822 707102 131004 707338
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 553254 120204 588698
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 373254 120204 408698
rect 119604 373018 119786 373254
rect 120022 373018 120204 373254
rect 119604 372934 120204 373018
rect 119604 372698 119786 372934
rect 120022 372698 120204 372934
rect 119604 337254 120204 372698
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7162 101786 -6926
rect 102022 -7162 102204 -6926
rect 101604 -7246 102204 -7162
rect 101604 -7482 101786 -7246
rect 102022 -7482 102204 -7246
rect 101604 -7504 102204 -7482
rect 119604 -5986 120204 12698
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 130404 672054 131004 707102
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3166 131004 23498
rect 130404 -3402 130586 -3166
rect 130822 -3402 131004 -3166
rect 130404 -3486 131004 -3402
rect 130404 -3722 130586 -3486
rect 130822 -3722 131004 -3486
rect 130404 -3744 131004 -3722
rect 134004 675654 134604 708982
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -5046 134604 27098
rect 134004 -5282 134186 -5046
rect 134422 -5282 134604 -5046
rect 134004 -5366 134604 -5282
rect 134004 -5602 134186 -5366
rect 134422 -5602 134604 -5366
rect 134004 -5624 134604 -5602
rect 137604 679254 138204 710862
rect 155604 710478 156204 711440
rect 155604 710242 155786 710478
rect 156022 710242 156204 710478
rect 155604 710158 156204 710242
rect 155604 709922 155786 710158
rect 156022 709922 156204 710158
rect 152004 708598 152604 709560
rect 152004 708362 152186 708598
rect 152422 708362 152604 708598
rect 152004 708278 152604 708362
rect 152004 708042 152186 708278
rect 152422 708042 152604 708278
rect 148404 706718 149004 707680
rect 148404 706482 148586 706718
rect 148822 706482 149004 706718
rect 148404 706398 149004 706482
rect 148404 706162 148586 706398
rect 148822 706162 149004 706398
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 535254 138204 570698
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6222 119786 -5986
rect 120022 -6222 120204 -5986
rect 119604 -6306 120204 -6222
rect 119604 -6542 119786 -6306
rect 120022 -6542 120204 -6306
rect 119604 -7504 120204 -6542
rect 137604 -6926 138204 30698
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 148404 690054 149004 706162
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2226 149004 5498
rect 148404 -2462 148586 -2226
rect 148822 -2462 149004 -2226
rect 148404 -2546 149004 -2462
rect 148404 -2782 148586 -2546
rect 148822 -2782 149004 -2546
rect 148404 -3744 149004 -2782
rect 152004 693654 152604 708042
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 155604 697254 156204 709922
rect 173604 711418 174204 711440
rect 173604 711182 173786 711418
rect 174022 711182 174204 711418
rect 173604 711098 174204 711182
rect 173604 710862 173786 711098
rect 174022 710862 174204 711098
rect 170004 709538 170604 709560
rect 170004 709302 170186 709538
rect 170422 709302 170604 709538
rect 170004 709218 170604 709302
rect 170004 708982 170186 709218
rect 170422 708982 170604 709218
rect 166404 707658 167004 707680
rect 166404 707422 166586 707658
rect 166822 707422 167004 707658
rect 166404 707338 167004 707422
rect 166404 707102 166586 707338
rect 166822 707102 167004 707338
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 411802 156204 444698
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 411802 163404 415898
rect 166404 672054 167004 707102
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 411802 167004 419498
rect 170004 675654 170604 708982
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 411802 170604 423098
rect 173604 679254 174204 710862
rect 191604 710478 192204 711440
rect 191604 710242 191786 710478
rect 192022 710242 192204 710478
rect 191604 710158 192204 710242
rect 191604 709922 191786 710158
rect 192022 709922 192204 710158
rect 188004 708598 188604 709560
rect 188004 708362 188186 708598
rect 188422 708362 188604 708598
rect 188004 708278 188604 708362
rect 188004 708042 188186 708278
rect 188422 708042 188604 708278
rect 184404 706718 185004 707680
rect 184404 706482 184586 706718
rect 184822 706482 185004 706718
rect 184404 706398 185004 706482
rect 184404 706162 184586 706398
rect 184822 706162 185004 706398
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 411802 174204 426698
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 411802 181404 433898
rect 184404 690054 185004 706162
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 411802 185004 437498
rect 188004 693654 188604 708042
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 411802 188604 441098
rect 191604 697254 192204 709922
rect 209604 711418 210204 711440
rect 209604 711182 209786 711418
rect 210022 711182 210204 711418
rect 209604 711098 210204 711182
rect 209604 710862 209786 711098
rect 210022 710862 210204 711098
rect 206004 709538 206604 709560
rect 206004 709302 206186 709538
rect 206422 709302 206604 709538
rect 206004 709218 206604 709302
rect 206004 708982 206186 709218
rect 206422 708982 206604 709218
rect 202404 707658 203004 707680
rect 202404 707422 202586 707658
rect 202822 707422 203004 707658
rect 202404 707338 203004 707422
rect 202404 707102 202586 707338
rect 202822 707102 203004 707338
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 411802 192204 444698
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 411802 199404 415898
rect 202404 672054 203004 707102
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 528054 203004 563498
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 202404 492054 203004 527498
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 411802 203004 419498
rect 206004 675654 206604 708982
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 531654 206604 567098
rect 206004 531418 206186 531654
rect 206422 531418 206604 531654
rect 206004 531334 206604 531418
rect 206004 531098 206186 531334
rect 206422 531098 206604 531334
rect 206004 495654 206604 531098
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 411802 206604 423098
rect 209604 679254 210204 710862
rect 227604 710478 228204 711440
rect 227604 710242 227786 710478
rect 228022 710242 228204 710478
rect 227604 710158 228204 710242
rect 227604 709922 227786 710158
rect 228022 709922 228204 710158
rect 224004 708598 224604 709560
rect 224004 708362 224186 708598
rect 224422 708362 224604 708598
rect 224004 708278 224604 708362
rect 224004 708042 224186 708278
rect 224422 708042 224604 708278
rect 220404 706718 221004 707680
rect 220404 706482 220586 706718
rect 220822 706482 221004 706718
rect 220404 706398 221004 706482
rect 220404 706162 220586 706398
rect 220822 706162 221004 706398
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 535254 210204 570698
rect 209604 535018 209786 535254
rect 210022 535018 210204 535254
rect 209604 534934 210204 535018
rect 209604 534698 209786 534934
rect 210022 534698 210204 534934
rect 209604 499254 210204 534698
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 411802 210204 426698
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 506454 217404 541898
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 411802 217404 433898
rect 220404 690054 221004 706162
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 411802 221004 437498
rect 224004 693654 224604 708042
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 549654 224604 585098
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 411802 224604 441098
rect 227604 697254 228204 709922
rect 245604 711418 246204 711440
rect 245604 711182 245786 711418
rect 246022 711182 246204 711418
rect 245604 711098 246204 711182
rect 245604 710862 245786 711098
rect 246022 710862 246204 711098
rect 242004 709538 242604 709560
rect 242004 709302 242186 709538
rect 242422 709302 242604 709538
rect 242004 709218 242604 709302
rect 242004 708982 242186 709218
rect 242422 708982 242604 709218
rect 238404 707658 239004 707680
rect 238404 707422 238586 707658
rect 238822 707422 239004 707658
rect 238404 707338 239004 707422
rect 238404 707102 238586 707338
rect 238822 707102 239004 707338
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 553254 228204 588698
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 411802 228204 444698
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 234804 411802 235404 415898
rect 238404 672054 239004 707102
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 564054 239004 599498
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 420054 239004 455498
rect 238404 419818 238586 420054
rect 238822 419818 239004 420054
rect 238404 419734 239004 419818
rect 238404 419498 238586 419734
rect 238822 419498 239004 419734
rect 238404 411802 239004 419498
rect 242004 675654 242604 708982
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 567654 242604 603098
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 242004 495654 242604 531098
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 242004 423654 242604 459098
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 242004 411802 242604 423098
rect 245604 679254 246204 710862
rect 263604 710478 264204 711440
rect 263604 710242 263786 710478
rect 264022 710242 264204 710478
rect 263604 710158 264204 710242
rect 263604 709922 263786 710158
rect 264022 709922 264204 710158
rect 260004 708598 260604 709560
rect 260004 708362 260186 708598
rect 260422 708362 260604 708598
rect 260004 708278 260604 708362
rect 260004 708042 260186 708278
rect 260422 708042 260604 708278
rect 256404 706718 257004 707680
rect 256404 706482 256586 706718
rect 256822 706482 257004 706718
rect 256404 706398 257004 706482
rect 256404 706162 256586 706398
rect 256822 706162 257004 706398
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 571254 246204 606698
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 535254 246204 570698
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 245604 499254 246204 534698
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 245604 427254 246204 462698
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 245604 411802 246204 426698
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 252804 411802 253404 433898
rect 256404 690054 257004 706162
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 411802 257004 437498
rect 260004 693654 260604 708042
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 477654 260604 513098
rect 260004 477418 260186 477654
rect 260422 477418 260604 477654
rect 260004 477334 260604 477418
rect 260004 477098 260186 477334
rect 260422 477098 260604 477334
rect 260004 441654 260604 477098
rect 260004 441418 260186 441654
rect 260422 441418 260604 441654
rect 260004 441334 260604 441418
rect 260004 441098 260186 441334
rect 260422 441098 260604 441334
rect 260004 411802 260604 441098
rect 263604 697254 264204 709922
rect 281604 711418 282204 711440
rect 281604 711182 281786 711418
rect 282022 711182 282204 711418
rect 281604 711098 282204 711182
rect 281604 710862 281786 711098
rect 282022 710862 282204 711098
rect 278004 709538 278604 709560
rect 278004 709302 278186 709538
rect 278422 709302 278604 709538
rect 278004 709218 278604 709302
rect 278004 708982 278186 709218
rect 278422 708982 278604 709218
rect 274404 707658 275004 707680
rect 274404 707422 274586 707658
rect 274822 707422 275004 707658
rect 274404 707338 275004 707422
rect 274404 707102 274586 707338
rect 274822 707102 275004 707338
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 517254 264204 552698
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 481254 264204 516698
rect 263604 481018 263786 481254
rect 264022 481018 264204 481254
rect 263604 480934 264204 481018
rect 263604 480698 263786 480934
rect 264022 480698 264204 480934
rect 263604 445254 264204 480698
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 411802 264204 444698
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 270804 411802 271404 415898
rect 274404 672054 275004 707102
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 420054 275004 455498
rect 274404 419818 274586 420054
rect 274822 419818 275004 420054
rect 274404 419734 275004 419818
rect 274404 419498 274586 419734
rect 274822 419498 275004 419734
rect 274404 411802 275004 419498
rect 278004 675654 278604 708982
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 459654 278604 495098
rect 278004 459418 278186 459654
rect 278422 459418 278604 459654
rect 278004 459334 278604 459418
rect 278004 459098 278186 459334
rect 278422 459098 278604 459334
rect 278004 423654 278604 459098
rect 278004 423418 278186 423654
rect 278422 423418 278604 423654
rect 278004 423334 278604 423418
rect 278004 423098 278186 423334
rect 278422 423098 278604 423334
rect 278004 411802 278604 423098
rect 281604 679254 282204 710862
rect 299604 710478 300204 711440
rect 299604 710242 299786 710478
rect 300022 710242 300204 710478
rect 299604 710158 300204 710242
rect 299604 709922 299786 710158
rect 300022 709922 300204 710158
rect 296004 708598 296604 709560
rect 296004 708362 296186 708598
rect 296422 708362 296604 708598
rect 296004 708278 296604 708362
rect 296004 708042 296186 708278
rect 296422 708042 296604 708278
rect 292404 706718 293004 707680
rect 292404 706482 292586 706718
rect 292822 706482 293004 706718
rect 292404 706398 293004 706482
rect 292404 706162 292586 706398
rect 292822 706162 293004 706398
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 463254 282204 498698
rect 281604 463018 281786 463254
rect 282022 463018 282204 463254
rect 281604 462934 282204 463018
rect 281604 462698 281786 462934
rect 282022 462698 282204 462934
rect 281604 427254 282204 462698
rect 281604 427018 281786 427254
rect 282022 427018 282204 427254
rect 281604 426934 282204 427018
rect 281604 426698 281786 426934
rect 282022 426698 282204 426934
rect 281604 411802 282204 426698
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 411802 289404 433898
rect 292404 690054 293004 706162
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 411802 293004 437498
rect 296004 693654 296604 708042
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 411802 296604 441098
rect 299604 697254 300204 709922
rect 317604 711418 318204 711440
rect 317604 711182 317786 711418
rect 318022 711182 318204 711418
rect 317604 711098 318204 711182
rect 317604 710862 317786 711098
rect 318022 710862 318204 711098
rect 314004 709538 314604 709560
rect 314004 709302 314186 709538
rect 314422 709302 314604 709538
rect 314004 709218 314604 709302
rect 314004 708982 314186 709218
rect 314422 708982 314604 709218
rect 310404 707658 311004 707680
rect 310404 707422 310586 707658
rect 310822 707422 311004 707658
rect 310404 707338 311004 707422
rect 310404 707102 310586 707338
rect 310822 707102 311004 707338
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 411802 300204 444698
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 411802 307404 415898
rect 310404 672054 311004 707102
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 310404 528054 311004 563498
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 411802 311004 419498
rect 314004 675654 314604 708982
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 567654 314604 603098
rect 314004 567418 314186 567654
rect 314422 567418 314604 567654
rect 314004 567334 314604 567418
rect 314004 567098 314186 567334
rect 314422 567098 314604 567334
rect 314004 531654 314604 567098
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 411802 314604 423098
rect 317604 679254 318204 710862
rect 335604 710478 336204 711440
rect 335604 710242 335786 710478
rect 336022 710242 336204 710478
rect 335604 710158 336204 710242
rect 335604 709922 335786 710158
rect 336022 709922 336204 710158
rect 332004 708598 332604 709560
rect 332004 708362 332186 708598
rect 332422 708362 332604 708598
rect 332004 708278 332604 708362
rect 332004 708042 332186 708278
rect 332422 708042 332604 708278
rect 328404 706718 329004 707680
rect 328404 706482 328586 706718
rect 328822 706482 329004 706718
rect 328404 706398 329004 706482
rect 328404 706162 328586 706398
rect 328822 706162 329004 706398
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 571254 318204 606698
rect 317604 571018 317786 571254
rect 318022 571018 318204 571254
rect 317604 570934 318204 571018
rect 317604 570698 317786 570934
rect 318022 570698 318204 570934
rect 317604 535254 318204 570698
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 411802 318204 426698
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 542454 325404 577898
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 411802 325404 433898
rect 328404 690054 329004 706162
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 546054 329004 581498
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 411802 329004 437498
rect 332004 693654 332604 708042
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 549654 332604 585098
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 513654 332604 549098
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 477654 332604 513098
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 411802 332604 441098
rect 335604 697254 336204 709922
rect 353604 711418 354204 711440
rect 353604 711182 353786 711418
rect 354022 711182 354204 711418
rect 353604 711098 354204 711182
rect 353604 710862 353786 711098
rect 354022 710862 354204 711098
rect 350004 709538 350604 709560
rect 350004 709302 350186 709538
rect 350422 709302 350604 709538
rect 350004 709218 350604 709302
rect 350004 708982 350186 709218
rect 350422 708982 350604 709218
rect 346404 707658 347004 707680
rect 346404 707422 346586 707658
rect 346822 707422 347004 707658
rect 346404 707338 347004 707422
rect 346404 707102 346586 707338
rect 346822 707102 347004 707338
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 553254 336204 588698
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 517254 336204 552698
rect 335604 517018 335786 517254
rect 336022 517018 336204 517254
rect 335604 516934 336204 517018
rect 335604 516698 335786 516934
rect 336022 516698 336204 516934
rect 335604 481254 336204 516698
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 411802 336204 444698
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 411802 343404 415898
rect 346404 672054 347004 707102
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 528054 347004 563498
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 411802 347004 419498
rect 350004 675654 350604 708982
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 567654 350604 603098
rect 350004 567418 350186 567654
rect 350422 567418 350604 567654
rect 350004 567334 350604 567418
rect 350004 567098 350186 567334
rect 350422 567098 350604 567334
rect 350004 531654 350604 567098
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 495654 350604 531098
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 411802 350604 423098
rect 353604 679254 354204 710862
rect 371604 710478 372204 711440
rect 371604 710242 371786 710478
rect 372022 710242 372204 710478
rect 371604 710158 372204 710242
rect 371604 709922 371786 710158
rect 372022 709922 372204 710158
rect 368004 708598 368604 709560
rect 368004 708362 368186 708598
rect 368422 708362 368604 708598
rect 368004 708278 368604 708362
rect 368004 708042 368186 708278
rect 368422 708042 368604 708278
rect 364404 706718 365004 707680
rect 364404 706482 364586 706718
rect 364822 706482 365004 706718
rect 364404 706398 365004 706482
rect 364404 706162 364586 706398
rect 364822 706162 365004 706398
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 571254 354204 606698
rect 353604 571018 353786 571254
rect 354022 571018 354204 571254
rect 353604 570934 354204 571018
rect 353604 570698 353786 570934
rect 354022 570698 354204 570934
rect 353604 535254 354204 570698
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 499254 354204 534698
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 411802 354204 426698
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 411802 361404 433898
rect 364404 690054 365004 706162
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 546054 365004 581498
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 510054 365004 545498
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 411802 365004 437498
rect 368004 693654 368604 708042
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 549654 368604 585098
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 513654 368604 549098
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 477654 368604 513098
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 411802 368604 441098
rect 371604 697254 372204 709922
rect 389604 711418 390204 711440
rect 389604 711182 389786 711418
rect 390022 711182 390204 711418
rect 389604 711098 390204 711182
rect 389604 710862 389786 711098
rect 390022 710862 390204 711098
rect 386004 709538 386604 709560
rect 386004 709302 386186 709538
rect 386422 709302 386604 709538
rect 386004 709218 386604 709302
rect 386004 708982 386186 709218
rect 386422 708982 386604 709218
rect 382404 707658 383004 707680
rect 382404 707422 382586 707658
rect 382822 707422 383004 707658
rect 382404 707338 383004 707422
rect 382404 707102 382586 707338
rect 382822 707102 383004 707338
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 553254 372204 588698
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 517254 372204 552698
rect 371604 517018 371786 517254
rect 372022 517018 372204 517254
rect 371604 516934 372204 517018
rect 371604 516698 371786 516934
rect 372022 516698 372204 516934
rect 371604 481254 372204 516698
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 411802 372204 444698
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 411802 379404 415898
rect 382404 672054 383004 707102
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 411802 383004 419498
rect 386004 675654 386604 708982
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 411802 386604 423098
rect 389604 679254 390204 710862
rect 407604 710478 408204 711440
rect 407604 710242 407786 710478
rect 408022 710242 408204 710478
rect 407604 710158 408204 710242
rect 407604 709922 407786 710158
rect 408022 709922 408204 710158
rect 404004 708598 404604 709560
rect 404004 708362 404186 708598
rect 404422 708362 404604 708598
rect 404004 708278 404604 708362
rect 404004 708042 404186 708278
rect 404422 708042 404604 708278
rect 400404 706718 401004 707680
rect 400404 706482 400586 706718
rect 400822 706482 401004 706718
rect 400404 706398 401004 706482
rect 400404 706162 400586 706398
rect 400822 706162 401004 706398
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 411802 390204 426698
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4106 152604 9098
rect 152004 -4342 152186 -4106
rect 152422 -4342 152604 -4106
rect 152004 -4426 152604 -4342
rect 152004 -4662 152186 -4426
rect 152422 -4662 152604 -4426
rect 152004 -5624 152604 -4662
rect 155604 157254 156204 175000
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7162 137786 -6926
rect 138022 -7162 138204 -6926
rect 137604 -7246 138204 -7162
rect 137604 -7482 137786 -7246
rect 138022 -7482 138204 -7246
rect 137604 -7504 138204 -7482
rect 155604 -5986 156204 12698
rect 162804 164454 163404 175000
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 166404 168054 167004 175000
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3166 167004 23498
rect 166404 -3402 166586 -3166
rect 166822 -3402 167004 -3166
rect 166404 -3486 167004 -3402
rect 166404 -3722 166586 -3486
rect 166822 -3722 167004 -3486
rect 166404 -3744 167004 -3722
rect 170004 171654 170604 175000
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -5046 170604 27098
rect 170004 -5282 170186 -5046
rect 170422 -5282 170604 -5046
rect 170004 -5366 170604 -5282
rect 170004 -5602 170186 -5366
rect 170422 -5602 170604 -5366
rect 170004 -5624 170604 -5602
rect 173604 139254 174204 175000
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6222 155786 -5986
rect 156022 -6222 156204 -5986
rect 155604 -6306 156204 -6222
rect 155604 -6542 155786 -6306
rect 156022 -6542 156204 -6306
rect 155604 -7504 156204 -6542
rect 173604 -6926 174204 30698
rect 180804 146454 181404 175000
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 184404 150054 185004 175000
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2226 185004 5498
rect 184404 -2462 184586 -2226
rect 184822 -2462 185004 -2226
rect 184404 -2546 185004 -2462
rect 184404 -2782 184586 -2546
rect 184822 -2782 185004 -2546
rect 184404 -3744 185004 -2782
rect 188004 153654 188604 175000
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4106 188604 9098
rect 188004 -4342 188186 -4106
rect 188422 -4342 188604 -4106
rect 188004 -4426 188604 -4342
rect 188004 -4662 188186 -4426
rect 188422 -4662 188604 -4426
rect 188004 -5624 188604 -4662
rect 191604 157254 192204 175000
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7162 173786 -6926
rect 174022 -7162 174204 -6926
rect 173604 -7246 174204 -7162
rect 173604 -7482 173786 -7246
rect 174022 -7482 174204 -7246
rect 173604 -7504 174204 -7482
rect 191604 -5986 192204 12698
rect 198804 164454 199404 175000
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 202404 168054 203004 175000
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3166 203004 23498
rect 202404 -3402 202586 -3166
rect 202822 -3402 203004 -3166
rect 202404 -3486 203004 -3402
rect 202404 -3722 202586 -3486
rect 202822 -3722 203004 -3486
rect 202404 -3744 203004 -3722
rect 206004 171654 206604 175000
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -5046 206604 27098
rect 206004 -5282 206186 -5046
rect 206422 -5282 206604 -5046
rect 206004 -5366 206604 -5282
rect 206004 -5602 206186 -5366
rect 206422 -5602 206604 -5366
rect 206004 -5624 206604 -5602
rect 209604 139254 210204 175000
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6222 191786 -5986
rect 192022 -6222 192204 -5986
rect 191604 -6306 192204 -6222
rect 191604 -6542 191786 -6306
rect 192022 -6542 192204 -6306
rect 191604 -7504 192204 -6542
rect 209604 -6926 210204 30698
rect 216804 146454 217404 175000
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 220404 150054 221004 175000
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2226 221004 5498
rect 220404 -2462 220586 -2226
rect 220822 -2462 221004 -2226
rect 220404 -2546 221004 -2462
rect 220404 -2782 220586 -2546
rect 220822 -2782 221004 -2546
rect 220404 -3744 221004 -2782
rect 224004 153654 224604 175000
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4106 224604 9098
rect 224004 -4342 224186 -4106
rect 224422 -4342 224604 -4106
rect 224004 -4426 224604 -4342
rect 224004 -4662 224186 -4426
rect 224422 -4662 224604 -4426
rect 224004 -5624 224604 -4662
rect 227604 157254 228204 175000
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7162 209786 -6926
rect 210022 -7162 210204 -6926
rect 209604 -7246 210204 -7162
rect 209604 -7482 209786 -7246
rect 210022 -7482 210204 -7246
rect 209604 -7504 210204 -7482
rect 227604 -5986 228204 12698
rect 234804 164454 235404 175000
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 238404 168054 239004 175000
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3166 239004 23498
rect 238404 -3402 238586 -3166
rect 238822 -3402 239004 -3166
rect 238404 -3486 239004 -3402
rect 238404 -3722 238586 -3486
rect 238822 -3722 239004 -3486
rect 238404 -3744 239004 -3722
rect 242004 171654 242604 175000
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -5046 242604 27098
rect 242004 -5282 242186 -5046
rect 242422 -5282 242604 -5046
rect 242004 -5366 242604 -5282
rect 242004 -5602 242186 -5366
rect 242422 -5602 242604 -5366
rect 242004 -5624 242604 -5602
rect 245604 139254 246204 175000
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6222 227786 -5986
rect 228022 -6222 228204 -5986
rect 227604 -6306 228204 -6222
rect 227604 -6542 227786 -6306
rect 228022 -6542 228204 -6306
rect 227604 -7504 228204 -6542
rect 245604 -6926 246204 30698
rect 252804 146454 253404 175000
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 256404 150054 257004 175000
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2226 257004 5498
rect 256404 -2462 256586 -2226
rect 256822 -2462 257004 -2226
rect 256404 -2546 257004 -2462
rect 256404 -2782 256586 -2546
rect 256822 -2782 257004 -2546
rect 256404 -3744 257004 -2782
rect 260004 153654 260604 175000
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4106 260604 9098
rect 260004 -4342 260186 -4106
rect 260422 -4342 260604 -4106
rect 260004 -4426 260604 -4342
rect 260004 -4662 260186 -4426
rect 260422 -4662 260604 -4426
rect 260004 -5624 260604 -4662
rect 263604 157254 264204 175000
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7162 245786 -6926
rect 246022 -7162 246204 -6926
rect 245604 -7246 246204 -7162
rect 245604 -7482 245786 -7246
rect 246022 -7482 246204 -7246
rect 245604 -7504 246204 -7482
rect 263604 -5986 264204 12698
rect 270804 164454 271404 175000
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 274404 168054 275004 175000
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3166 275004 23498
rect 274404 -3402 274586 -3166
rect 274822 -3402 275004 -3166
rect 274404 -3486 275004 -3402
rect 274404 -3722 274586 -3486
rect 274822 -3722 275004 -3486
rect 274404 -3744 275004 -3722
rect 278004 171654 278604 175000
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -5046 278604 27098
rect 278004 -5282 278186 -5046
rect 278422 -5282 278604 -5046
rect 278004 -5366 278604 -5282
rect 278004 -5602 278186 -5366
rect 278422 -5602 278604 -5366
rect 278004 -5624 278604 -5602
rect 281604 139254 282204 175000
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6222 263786 -5986
rect 264022 -6222 264204 -5986
rect 263604 -6306 264204 -6222
rect 263604 -6542 263786 -6306
rect 264022 -6542 264204 -6306
rect 263604 -7504 264204 -6542
rect 281604 -6926 282204 30698
rect 288804 146454 289404 175000
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 292404 150054 293004 175000
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2226 293004 5498
rect 292404 -2462 292586 -2226
rect 292822 -2462 293004 -2226
rect 292404 -2546 293004 -2462
rect 292404 -2782 292586 -2546
rect 292822 -2782 293004 -2546
rect 292404 -3744 293004 -2782
rect 296004 153654 296604 175000
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4106 296604 9098
rect 296004 -4342 296186 -4106
rect 296422 -4342 296604 -4106
rect 296004 -4426 296604 -4342
rect 296004 -4662 296186 -4426
rect 296422 -4662 296604 -4426
rect 296004 -5624 296604 -4662
rect 299604 157254 300204 175000
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7162 281786 -6926
rect 282022 -7162 282204 -6926
rect 281604 -7246 282204 -7162
rect 281604 -7482 281786 -7246
rect 282022 -7482 282204 -7246
rect 281604 -7504 282204 -7482
rect 299604 -5986 300204 12698
rect 306804 164454 307404 175000
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 310404 168054 311004 175000
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3166 311004 23498
rect 310404 -3402 310586 -3166
rect 310822 -3402 311004 -3166
rect 310404 -3486 311004 -3402
rect 310404 -3722 310586 -3486
rect 310822 -3722 311004 -3486
rect 310404 -3744 311004 -3722
rect 314004 171654 314604 175000
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -5046 314604 27098
rect 314004 -5282 314186 -5046
rect 314422 -5282 314604 -5046
rect 314004 -5366 314604 -5282
rect 314004 -5602 314186 -5366
rect 314422 -5602 314604 -5366
rect 314004 -5624 314604 -5602
rect 317604 139254 318204 175000
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 317604 103254 318204 138698
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6222 299786 -5986
rect 300022 -6222 300204 -5986
rect 299604 -6306 300204 -6222
rect 299604 -6542 299786 -6306
rect 300022 -6542 300204 -6306
rect 299604 -7504 300204 -6542
rect 317604 -6926 318204 30698
rect 324804 146454 325404 175000
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 328404 150054 329004 175000
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2226 329004 5498
rect 328404 -2462 328586 -2226
rect 328822 -2462 329004 -2226
rect 328404 -2546 329004 -2462
rect 328404 -2782 328586 -2546
rect 328822 -2782 329004 -2546
rect 328404 -3744 329004 -2782
rect 332004 153654 332604 175000
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 332004 117654 332604 153098
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4106 332604 9098
rect 332004 -4342 332186 -4106
rect 332422 -4342 332604 -4106
rect 332004 -4426 332604 -4342
rect 332004 -4662 332186 -4426
rect 332422 -4662 332604 -4426
rect 332004 -5624 332604 -4662
rect 335604 157254 336204 175000
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7162 317786 -6926
rect 318022 -7162 318204 -6926
rect 317604 -7246 318204 -7162
rect 317604 -7482 317786 -7246
rect 318022 -7482 318204 -7246
rect 317604 -7504 318204 -7482
rect 335604 -5986 336204 12698
rect 342804 164454 343404 175000
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 346404 168054 347004 175000
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3166 347004 23498
rect 346404 -3402 346586 -3166
rect 346822 -3402 347004 -3166
rect 346404 -3486 347004 -3402
rect 346404 -3722 346586 -3486
rect 346822 -3722 347004 -3486
rect 346404 -3744 347004 -3722
rect 350004 171654 350604 175000
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -5046 350604 27098
rect 350004 -5282 350186 -5046
rect 350422 -5282 350604 -5046
rect 350004 -5366 350604 -5282
rect 350004 -5602 350186 -5366
rect 350422 -5602 350604 -5366
rect 350004 -5624 350604 -5602
rect 353604 139254 354204 175000
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6222 335786 -5986
rect 336022 -6222 336204 -5986
rect 335604 -6306 336204 -6222
rect 335604 -6542 335786 -6306
rect 336022 -6542 336204 -6306
rect 335604 -7504 336204 -6542
rect 353604 -6926 354204 30698
rect 360804 146454 361404 175000
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 364404 150054 365004 175000
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2226 365004 5498
rect 364404 -2462 364586 -2226
rect 364822 -2462 365004 -2226
rect 364404 -2546 365004 -2462
rect 364404 -2782 364586 -2546
rect 364822 -2782 365004 -2546
rect 364404 -3744 365004 -2782
rect 368004 153654 368604 175000
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 368004 117654 368604 153098
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4106 368604 9098
rect 368004 -4342 368186 -4106
rect 368422 -4342 368604 -4106
rect 368004 -4426 368604 -4342
rect 368004 -4662 368186 -4426
rect 368422 -4662 368604 -4426
rect 368004 -5624 368604 -4662
rect 371604 157254 372204 175000
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 371604 121254 372204 156698
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7162 353786 -6926
rect 354022 -7162 354204 -6926
rect 353604 -7246 354204 -7162
rect 353604 -7482 353786 -7246
rect 354022 -7482 354204 -7246
rect 353604 -7504 354204 -7482
rect 371604 -5986 372204 12698
rect 378804 164454 379404 175000
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 382404 168054 383004 175000
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 386004 171654 386604 175000
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 384987 66196 385053 66197
rect 384987 66132 384988 66196
rect 385052 66132 385053 66196
rect 384987 66131 385053 66132
rect 384990 60621 385050 66131
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 384987 60620 385053 60621
rect 384987 60556 384988 60620
rect 385052 60556 385053 60620
rect 384987 60555 385053 60556
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3166 383004 23498
rect 382404 -3402 382586 -3166
rect 382822 -3402 383004 -3166
rect 382404 -3486 383004 -3402
rect 382404 -3722 382586 -3486
rect 382822 -3722 383004 -3486
rect 382404 -3744 383004 -3722
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -5046 386604 27098
rect 386004 -5282 386186 -5046
rect 386422 -5282 386604 -5046
rect 386004 -5366 386604 -5282
rect 386004 -5602 386186 -5366
rect 386422 -5602 386604 -5366
rect 386004 -5624 386604 -5602
rect 389604 139254 390204 175000
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6222 371786 -5986
rect 372022 -6222 372204 -5986
rect 371604 -6306 372204 -6222
rect 371604 -6542 371786 -6306
rect 372022 -6542 372204 -6306
rect 371604 -7504 372204 -6542
rect 389604 -6926 390204 30698
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 400404 690054 401004 706162
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 366054 401004 401498
rect 400404 365818 400586 366054
rect 400822 365818 401004 366054
rect 400404 365734 401004 365818
rect 400404 365498 400586 365734
rect 400822 365498 401004 365734
rect 400404 330054 401004 365498
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2226 401004 5498
rect 400404 -2462 400586 -2226
rect 400822 -2462 401004 -2226
rect 400404 -2546 401004 -2462
rect 400404 -2782 400586 -2546
rect 400822 -2782 401004 -2546
rect 400404 -3744 401004 -2782
rect 404004 693654 404604 708042
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 369654 404604 405098
rect 404004 369418 404186 369654
rect 404422 369418 404604 369654
rect 404004 369334 404604 369418
rect 404004 369098 404186 369334
rect 404422 369098 404604 369334
rect 404004 333654 404604 369098
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 297654 404604 333098
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4106 404604 9098
rect 404004 -4342 404186 -4106
rect 404422 -4342 404604 -4106
rect 404004 -4426 404604 -4342
rect 404004 -4662 404186 -4426
rect 404422 -4662 404604 -4426
rect 404004 -5624 404604 -4662
rect 407604 697254 408204 709922
rect 425604 711418 426204 711440
rect 425604 711182 425786 711418
rect 426022 711182 426204 711418
rect 425604 711098 426204 711182
rect 425604 710862 425786 711098
rect 426022 710862 426204 711098
rect 422004 709538 422604 709560
rect 422004 709302 422186 709538
rect 422422 709302 422604 709538
rect 422004 709218 422604 709302
rect 422004 708982 422186 709218
rect 422422 708982 422604 709218
rect 418404 707658 419004 707680
rect 418404 707422 418586 707658
rect 418822 707422 419004 707658
rect 418404 707338 419004 707422
rect 418404 707102 418586 707338
rect 418822 707102 419004 707338
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 373254 408204 408698
rect 407604 373018 407786 373254
rect 408022 373018 408204 373254
rect 407604 372934 408204 373018
rect 407604 372698 407786 372934
rect 408022 372698 408204 372934
rect 407604 337254 408204 372698
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 301254 408204 336698
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7162 389786 -6926
rect 390022 -7162 390204 -6926
rect 389604 -7246 390204 -7162
rect 389604 -7482 389786 -7246
rect 390022 -7482 390204 -7246
rect 389604 -7504 390204 -7482
rect 407604 -5986 408204 12698
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 418404 672054 419004 707102
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3166 419004 23498
rect 418404 -3402 418586 -3166
rect 418822 -3402 419004 -3166
rect 418404 -3486 419004 -3402
rect 418404 -3722 418586 -3486
rect 418822 -3722 419004 -3486
rect 418404 -3744 419004 -3722
rect 422004 675654 422604 708982
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -5046 422604 27098
rect 422004 -5282 422186 -5046
rect 422422 -5282 422604 -5046
rect 422004 -5366 422604 -5282
rect 422004 -5602 422186 -5366
rect 422422 -5602 422604 -5366
rect 422004 -5624 422604 -5602
rect 425604 679254 426204 710862
rect 443604 710478 444204 711440
rect 443604 710242 443786 710478
rect 444022 710242 444204 710478
rect 443604 710158 444204 710242
rect 443604 709922 443786 710158
rect 444022 709922 444204 710158
rect 440004 708598 440604 709560
rect 440004 708362 440186 708598
rect 440422 708362 440604 708598
rect 440004 708278 440604 708362
rect 440004 708042 440186 708278
rect 440422 708042 440604 708278
rect 436404 706718 437004 707680
rect 436404 706482 436586 706718
rect 436822 706482 437004 706718
rect 436404 706398 437004 706482
rect 436404 706162 436586 706398
rect 436822 706162 437004 706398
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6222 407786 -5986
rect 408022 -6222 408204 -5986
rect 407604 -6306 408204 -6222
rect 407604 -6542 407786 -6306
rect 408022 -6542 408204 -6306
rect 407604 -7504 408204 -6542
rect 425604 -6926 426204 30698
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 436404 690054 437004 706162
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2226 437004 5498
rect 436404 -2462 436586 -2226
rect 436822 -2462 437004 -2226
rect 436404 -2546 437004 -2462
rect 436404 -2782 436586 -2546
rect 436822 -2782 437004 -2546
rect 436404 -3744 437004 -2782
rect 440004 693654 440604 708042
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4106 440604 9098
rect 440004 -4342 440186 -4106
rect 440422 -4342 440604 -4106
rect 440004 -4426 440604 -4342
rect 440004 -4662 440186 -4426
rect 440422 -4662 440604 -4426
rect 440004 -5624 440604 -4662
rect 443604 697254 444204 709922
rect 461604 711418 462204 711440
rect 461604 711182 461786 711418
rect 462022 711182 462204 711418
rect 461604 711098 462204 711182
rect 461604 710862 461786 711098
rect 462022 710862 462204 711098
rect 458004 709538 458604 709560
rect 458004 709302 458186 709538
rect 458422 709302 458604 709538
rect 458004 709218 458604 709302
rect 458004 708982 458186 709218
rect 458422 708982 458604 709218
rect 454404 707658 455004 707680
rect 454404 707422 454586 707658
rect 454822 707422 455004 707658
rect 454404 707338 455004 707422
rect 454404 707102 454586 707338
rect 454822 707102 455004 707338
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7162 425786 -6926
rect 426022 -7162 426204 -6926
rect 425604 -7246 426204 -7162
rect 425604 -7482 425786 -7246
rect 426022 -7482 426204 -7246
rect 425604 -7504 426204 -7482
rect 443604 -5986 444204 12698
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 454404 672054 455004 707102
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3166 455004 23498
rect 454404 -3402 454586 -3166
rect 454822 -3402 455004 -3166
rect 454404 -3486 455004 -3402
rect 454404 -3722 454586 -3486
rect 454822 -3722 455004 -3486
rect 454404 -3744 455004 -3722
rect 458004 675654 458604 708982
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -5046 458604 27098
rect 458004 -5282 458186 -5046
rect 458422 -5282 458604 -5046
rect 458004 -5366 458604 -5282
rect 458004 -5602 458186 -5366
rect 458422 -5602 458604 -5366
rect 458004 -5624 458604 -5602
rect 461604 679254 462204 710862
rect 479604 710478 480204 711440
rect 479604 710242 479786 710478
rect 480022 710242 480204 710478
rect 479604 710158 480204 710242
rect 479604 709922 479786 710158
rect 480022 709922 480204 710158
rect 476004 708598 476604 709560
rect 476004 708362 476186 708598
rect 476422 708362 476604 708598
rect 476004 708278 476604 708362
rect 476004 708042 476186 708278
rect 476422 708042 476604 708278
rect 472404 706718 473004 707680
rect 472404 706482 472586 706718
rect 472822 706482 473004 706718
rect 472404 706398 473004 706482
rect 472404 706162 472586 706398
rect 472822 706162 473004 706398
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6222 443786 -5986
rect 444022 -6222 444204 -5986
rect 443604 -6306 444204 -6222
rect 443604 -6542 443786 -6306
rect 444022 -6542 444204 -6306
rect 443604 -7504 444204 -6542
rect 461604 -6926 462204 30698
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 472404 690054 473004 706162
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2226 473004 5498
rect 472404 -2462 472586 -2226
rect 472822 -2462 473004 -2226
rect 472404 -2546 473004 -2462
rect 472404 -2782 472586 -2546
rect 472822 -2782 473004 -2546
rect 472404 -3744 473004 -2782
rect 476004 693654 476604 708042
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4106 476604 9098
rect 476004 -4342 476186 -4106
rect 476422 -4342 476604 -4106
rect 476004 -4426 476604 -4342
rect 476004 -4662 476186 -4426
rect 476422 -4662 476604 -4426
rect 476004 -5624 476604 -4662
rect 479604 697254 480204 709922
rect 497604 711418 498204 711440
rect 497604 711182 497786 711418
rect 498022 711182 498204 711418
rect 497604 711098 498204 711182
rect 497604 710862 497786 711098
rect 498022 710862 498204 711098
rect 494004 709538 494604 709560
rect 494004 709302 494186 709538
rect 494422 709302 494604 709538
rect 494004 709218 494604 709302
rect 494004 708982 494186 709218
rect 494422 708982 494604 709218
rect 490404 707658 491004 707680
rect 490404 707422 490586 707658
rect 490822 707422 491004 707658
rect 490404 707338 491004 707422
rect 490404 707102 490586 707338
rect 490822 707102 491004 707338
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 553254 480204 588698
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7162 461786 -6926
rect 462022 -7162 462204 -6926
rect 461604 -7246 462204 -7162
rect 461604 -7482 461786 -7246
rect 462022 -7482 462204 -7246
rect 461604 -7504 462204 -7482
rect 479604 -5986 480204 12698
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 490404 672054 491004 707102
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3166 491004 23498
rect 490404 -3402 490586 -3166
rect 490822 -3402 491004 -3166
rect 490404 -3486 491004 -3402
rect 490404 -3722 490586 -3486
rect 490822 -3722 491004 -3486
rect 490404 -3744 491004 -3722
rect 494004 675654 494604 708982
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 531654 494604 567098
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -5046 494604 27098
rect 494004 -5282 494186 -5046
rect 494422 -5282 494604 -5046
rect 494004 -5366 494604 -5282
rect 494004 -5602 494186 -5366
rect 494422 -5602 494604 -5366
rect 494004 -5624 494604 -5602
rect 497604 679254 498204 710862
rect 515604 710478 516204 711440
rect 515604 710242 515786 710478
rect 516022 710242 516204 710478
rect 515604 710158 516204 710242
rect 515604 709922 515786 710158
rect 516022 709922 516204 710158
rect 512004 708598 512604 709560
rect 512004 708362 512186 708598
rect 512422 708362 512604 708598
rect 512004 708278 512604 708362
rect 512004 708042 512186 708278
rect 512422 708042 512604 708278
rect 508404 706718 509004 707680
rect 508404 706482 508586 706718
rect 508822 706482 509004 706718
rect 508404 706398 509004 706482
rect 508404 706162 508586 706398
rect 508822 706162 509004 706398
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 535254 498204 570698
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6222 479786 -5986
rect 480022 -6222 480204 -5986
rect 479604 -6306 480204 -6222
rect 479604 -6542 479786 -6306
rect 480022 -6542 480204 -6306
rect 479604 -7504 480204 -6542
rect 497604 -6926 498204 30698
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 508404 690054 509004 706162
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2226 509004 5498
rect 508404 -2462 508586 -2226
rect 508822 -2462 509004 -2226
rect 508404 -2546 509004 -2462
rect 508404 -2782 508586 -2546
rect 508822 -2782 509004 -2546
rect 508404 -3744 509004 -2782
rect 512004 693654 512604 708042
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4106 512604 9098
rect 512004 -4342 512186 -4106
rect 512422 -4342 512604 -4106
rect 512004 -4426 512604 -4342
rect 512004 -4662 512186 -4426
rect 512422 -4662 512604 -4426
rect 512004 -5624 512604 -4662
rect 515604 697254 516204 709922
rect 533604 711418 534204 711440
rect 533604 711182 533786 711418
rect 534022 711182 534204 711418
rect 533604 711098 534204 711182
rect 533604 710862 533786 711098
rect 534022 710862 534204 711098
rect 530004 709538 530604 709560
rect 530004 709302 530186 709538
rect 530422 709302 530604 709538
rect 530004 709218 530604 709302
rect 530004 708982 530186 709218
rect 530422 708982 530604 709218
rect 526404 707658 527004 707680
rect 526404 707422 526586 707658
rect 526822 707422 527004 707658
rect 526404 707338 527004 707422
rect 526404 707102 526586 707338
rect 526822 707102 527004 707338
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7162 497786 -6926
rect 498022 -7162 498204 -6926
rect 497604 -7246 498204 -7162
rect 497604 -7482 497786 -7246
rect 498022 -7482 498204 -7246
rect 497604 -7504 498204 -7482
rect 515604 -5986 516204 12698
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 526404 672054 527004 707102
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3166 527004 23498
rect 526404 -3402 526586 -3166
rect 526822 -3402 527004 -3166
rect 526404 -3486 527004 -3402
rect 526404 -3722 526586 -3486
rect 526822 -3722 527004 -3486
rect 526404 -3744 527004 -3722
rect 530004 675654 530604 708982
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -5046 530604 27098
rect 530004 -5282 530186 -5046
rect 530422 -5282 530604 -5046
rect 530004 -5366 530604 -5282
rect 530004 -5602 530186 -5366
rect 530422 -5602 530604 -5366
rect 530004 -5624 530604 -5602
rect 533604 679254 534204 710862
rect 551604 710478 552204 711440
rect 551604 710242 551786 710478
rect 552022 710242 552204 710478
rect 551604 710158 552204 710242
rect 551604 709922 551786 710158
rect 552022 709922 552204 710158
rect 548004 708598 548604 709560
rect 548004 708362 548186 708598
rect 548422 708362 548604 708598
rect 548004 708278 548604 708362
rect 548004 708042 548186 708278
rect 548422 708042 548604 708278
rect 544404 706718 545004 707680
rect 544404 706482 544586 706718
rect 544822 706482 545004 706718
rect 544404 706398 545004 706482
rect 544404 706162 544586 706398
rect 544822 706162 545004 706398
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6222 515786 -5986
rect 516022 -6222 516204 -5986
rect 515604 -6306 516204 -6222
rect 515604 -6542 515786 -6306
rect 516022 -6542 516204 -6306
rect 515604 -7504 516204 -6542
rect 533604 -6926 534204 30698
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 544404 690054 545004 706162
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2226 545004 5498
rect 544404 -2462 544586 -2226
rect 544822 -2462 545004 -2226
rect 544404 -2546 545004 -2462
rect 544404 -2782 544586 -2546
rect 544822 -2782 545004 -2546
rect 544404 -3744 545004 -2782
rect 548004 693654 548604 708042
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4106 548604 9098
rect 548004 -4342 548186 -4106
rect 548422 -4342 548604 -4106
rect 548004 -4426 548604 -4342
rect 548004 -4662 548186 -4426
rect 548422 -4662 548604 -4426
rect 548004 -5624 548604 -4662
rect 551604 697254 552204 709922
rect 569604 711418 570204 711440
rect 569604 711182 569786 711418
rect 570022 711182 570204 711418
rect 569604 711098 570204 711182
rect 569604 710862 569786 711098
rect 570022 710862 570204 711098
rect 566004 709538 566604 709560
rect 566004 709302 566186 709538
rect 566422 709302 566604 709538
rect 566004 709218 566604 709302
rect 566004 708982 566186 709218
rect 566422 708982 566604 709218
rect 562404 707658 563004 707680
rect 562404 707422 562586 707658
rect 562822 707422 563004 707658
rect 562404 707338 563004 707422
rect 562404 707102 562586 707338
rect 562822 707102 563004 707338
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7162 533786 -6926
rect 534022 -7162 534204 -6926
rect 533604 -7246 534204 -7162
rect 533604 -7482 533786 -7246
rect 534022 -7482 534204 -7246
rect 533604 -7504 534204 -7482
rect 551604 -5986 552204 12698
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 562404 672054 563004 707102
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3166 563004 23498
rect 562404 -3402 562586 -3166
rect 562822 -3402 563004 -3166
rect 562404 -3486 563004 -3402
rect 562404 -3722 562586 -3486
rect 562822 -3722 563004 -3486
rect 562404 -3744 563004 -3722
rect 566004 675654 566604 708982
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -5046 566604 27098
rect 566004 -5282 566186 -5046
rect 566422 -5282 566604 -5046
rect 566004 -5366 566604 -5282
rect 566004 -5602 566186 -5366
rect 566422 -5602 566604 -5366
rect 566004 -5624 566604 -5602
rect 569604 679254 570204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 580404 706718 581004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 580404 706482 580586 706718
rect 580822 706482 581004 706718
rect 580404 706398 581004 706482
rect 580404 706162 580586 706398
rect 580822 706162 581004 706398
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6222 551786 -5986
rect 552022 -6222 552204 -5986
rect 551604 -6306 552204 -6222
rect 551604 -6542 551786 -6306
rect 552022 -6542 552204 -6306
rect 551604 -7504 552204 -6542
rect 569604 -6926 570204 30698
rect 576804 704838 577404 705800
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 580404 690054 581004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2226 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 690054 587800 706162
rect 587200 689818 587382 690054
rect 587618 689818 587800 690054
rect 587200 689734 587800 689818
rect 587200 689498 587382 689734
rect 587618 689498 587800 689734
rect 587200 654054 587800 689498
rect 587200 653818 587382 654054
rect 587618 653818 587800 654054
rect 587200 653734 587800 653818
rect 587200 653498 587382 653734
rect 587618 653498 587800 653734
rect 587200 618054 587800 653498
rect 587200 617818 587382 618054
rect 587618 617818 587800 618054
rect 587200 617734 587800 617818
rect 587200 617498 587382 617734
rect 587618 617498 587800 617734
rect 587200 582054 587800 617498
rect 587200 581818 587382 582054
rect 587618 581818 587800 582054
rect 587200 581734 587800 581818
rect 587200 581498 587382 581734
rect 587618 581498 587800 581734
rect 587200 546054 587800 581498
rect 587200 545818 587382 546054
rect 587618 545818 587800 546054
rect 587200 545734 587800 545818
rect 587200 545498 587382 545734
rect 587618 545498 587800 545734
rect 587200 510054 587800 545498
rect 587200 509818 587382 510054
rect 587618 509818 587800 510054
rect 587200 509734 587800 509818
rect 587200 509498 587382 509734
rect 587618 509498 587800 509734
rect 587200 474054 587800 509498
rect 587200 473818 587382 474054
rect 587618 473818 587800 474054
rect 587200 473734 587800 473818
rect 587200 473498 587382 473734
rect 587618 473498 587800 473734
rect 587200 438054 587800 473498
rect 587200 437818 587382 438054
rect 587618 437818 587800 438054
rect 587200 437734 587800 437818
rect 587200 437498 587382 437734
rect 587618 437498 587800 437734
rect 587200 402054 587800 437498
rect 587200 401818 587382 402054
rect 587618 401818 587800 402054
rect 587200 401734 587800 401818
rect 587200 401498 587382 401734
rect 587618 401498 587800 401734
rect 587200 366054 587800 401498
rect 587200 365818 587382 366054
rect 587618 365818 587800 366054
rect 587200 365734 587800 365818
rect 587200 365498 587382 365734
rect 587618 365498 587800 365734
rect 587200 330054 587800 365498
rect 587200 329818 587382 330054
rect 587618 329818 587800 330054
rect 587200 329734 587800 329818
rect 587200 329498 587382 329734
rect 587618 329498 587800 329734
rect 587200 294054 587800 329498
rect 587200 293818 587382 294054
rect 587618 293818 587800 294054
rect 587200 293734 587800 293818
rect 587200 293498 587382 293734
rect 587618 293498 587800 293734
rect 587200 258054 587800 293498
rect 587200 257818 587382 258054
rect 587618 257818 587800 258054
rect 587200 257734 587800 257818
rect 587200 257498 587382 257734
rect 587618 257498 587800 257734
rect 587200 222054 587800 257498
rect 587200 221818 587382 222054
rect 587618 221818 587800 222054
rect 587200 221734 587800 221818
rect 587200 221498 587382 221734
rect 587618 221498 587800 221734
rect 587200 186054 587800 221498
rect 587200 185818 587382 186054
rect 587618 185818 587800 186054
rect 587200 185734 587800 185818
rect 587200 185498 587382 185734
rect 587618 185498 587800 185734
rect 587200 150054 587800 185498
rect 587200 149818 587382 150054
rect 587618 149818 587800 150054
rect 587200 149734 587800 149818
rect 587200 149498 587382 149734
rect 587618 149498 587800 149734
rect 587200 114054 587800 149498
rect 587200 113818 587382 114054
rect 587618 113818 587800 114054
rect 587200 113734 587800 113818
rect 587200 113498 587382 113734
rect 587618 113498 587800 113734
rect 587200 78054 587800 113498
rect 587200 77818 587382 78054
rect 587618 77818 587800 78054
rect 587200 77734 587800 77818
rect 587200 77498 587382 77734
rect 587618 77498 587800 77734
rect 587200 42054 587800 77498
rect 587200 41818 587382 42054
rect 587618 41818 587800 42054
rect 587200 41734 587800 41818
rect 587200 41498 587382 41734
rect 587618 41498 587800 41734
rect 587200 6054 587800 41498
rect 587200 5818 587382 6054
rect 587618 5818 587800 6054
rect 587200 5734 587800 5818
rect 587200 5498 587382 5734
rect 587618 5498 587800 5734
rect 580404 -2462 580586 -2226
rect 580822 -2462 581004 -2226
rect 580404 -2546 581004 -2462
rect 580404 -2782 580586 -2546
rect 580822 -2782 581004 -2546
rect 580404 -3744 581004 -2782
rect 587200 -2226 587800 5498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 672054 588740 707102
rect 588140 671818 588322 672054
rect 588558 671818 588740 672054
rect 588140 671734 588740 671818
rect 588140 671498 588322 671734
rect 588558 671498 588740 671734
rect 588140 636054 588740 671498
rect 588140 635818 588322 636054
rect 588558 635818 588740 636054
rect 588140 635734 588740 635818
rect 588140 635498 588322 635734
rect 588558 635498 588740 635734
rect 588140 600054 588740 635498
rect 588140 599818 588322 600054
rect 588558 599818 588740 600054
rect 588140 599734 588740 599818
rect 588140 599498 588322 599734
rect 588558 599498 588740 599734
rect 588140 564054 588740 599498
rect 588140 563818 588322 564054
rect 588558 563818 588740 564054
rect 588140 563734 588740 563818
rect 588140 563498 588322 563734
rect 588558 563498 588740 563734
rect 588140 528054 588740 563498
rect 588140 527818 588322 528054
rect 588558 527818 588740 528054
rect 588140 527734 588740 527818
rect 588140 527498 588322 527734
rect 588558 527498 588740 527734
rect 588140 492054 588740 527498
rect 588140 491818 588322 492054
rect 588558 491818 588740 492054
rect 588140 491734 588740 491818
rect 588140 491498 588322 491734
rect 588558 491498 588740 491734
rect 588140 456054 588740 491498
rect 588140 455818 588322 456054
rect 588558 455818 588740 456054
rect 588140 455734 588740 455818
rect 588140 455498 588322 455734
rect 588558 455498 588740 455734
rect 588140 420054 588740 455498
rect 588140 419818 588322 420054
rect 588558 419818 588740 420054
rect 588140 419734 588740 419818
rect 588140 419498 588322 419734
rect 588558 419498 588740 419734
rect 588140 384054 588740 419498
rect 588140 383818 588322 384054
rect 588558 383818 588740 384054
rect 588140 383734 588740 383818
rect 588140 383498 588322 383734
rect 588558 383498 588740 383734
rect 588140 348054 588740 383498
rect 588140 347818 588322 348054
rect 588558 347818 588740 348054
rect 588140 347734 588740 347818
rect 588140 347498 588322 347734
rect 588558 347498 588740 347734
rect 588140 312054 588740 347498
rect 588140 311818 588322 312054
rect 588558 311818 588740 312054
rect 588140 311734 588740 311818
rect 588140 311498 588322 311734
rect 588558 311498 588740 311734
rect 588140 276054 588740 311498
rect 588140 275818 588322 276054
rect 588558 275818 588740 276054
rect 588140 275734 588740 275818
rect 588140 275498 588322 275734
rect 588558 275498 588740 275734
rect 588140 240054 588740 275498
rect 588140 239818 588322 240054
rect 588558 239818 588740 240054
rect 588140 239734 588740 239818
rect 588140 239498 588322 239734
rect 588558 239498 588740 239734
rect 588140 204054 588740 239498
rect 588140 203818 588322 204054
rect 588558 203818 588740 204054
rect 588140 203734 588740 203818
rect 588140 203498 588322 203734
rect 588558 203498 588740 203734
rect 588140 168054 588740 203498
rect 588140 167818 588322 168054
rect 588558 167818 588740 168054
rect 588140 167734 588740 167818
rect 588140 167498 588322 167734
rect 588558 167498 588740 167734
rect 588140 132054 588740 167498
rect 588140 131818 588322 132054
rect 588558 131818 588740 132054
rect 588140 131734 588740 131818
rect 588140 131498 588322 131734
rect 588558 131498 588740 131734
rect 588140 96054 588740 131498
rect 588140 95818 588322 96054
rect 588558 95818 588740 96054
rect 588140 95734 588740 95818
rect 588140 95498 588322 95734
rect 588558 95498 588740 95734
rect 588140 60054 588740 95498
rect 588140 59818 588322 60054
rect 588558 59818 588740 60054
rect 588140 59734 588740 59818
rect 588140 59498 588322 59734
rect 588558 59498 588740 59734
rect 588140 24054 588740 59498
rect 588140 23818 588322 24054
rect 588558 23818 588740 24054
rect 588140 23734 588740 23818
rect 588140 23498 588322 23734
rect 588558 23498 588740 23734
rect 588140 -3166 588740 23498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 693654 589680 708042
rect 589080 693418 589262 693654
rect 589498 693418 589680 693654
rect 589080 693334 589680 693418
rect 589080 693098 589262 693334
rect 589498 693098 589680 693334
rect 589080 657654 589680 693098
rect 589080 657418 589262 657654
rect 589498 657418 589680 657654
rect 589080 657334 589680 657418
rect 589080 657098 589262 657334
rect 589498 657098 589680 657334
rect 589080 621654 589680 657098
rect 589080 621418 589262 621654
rect 589498 621418 589680 621654
rect 589080 621334 589680 621418
rect 589080 621098 589262 621334
rect 589498 621098 589680 621334
rect 589080 585654 589680 621098
rect 589080 585418 589262 585654
rect 589498 585418 589680 585654
rect 589080 585334 589680 585418
rect 589080 585098 589262 585334
rect 589498 585098 589680 585334
rect 589080 549654 589680 585098
rect 589080 549418 589262 549654
rect 589498 549418 589680 549654
rect 589080 549334 589680 549418
rect 589080 549098 589262 549334
rect 589498 549098 589680 549334
rect 589080 513654 589680 549098
rect 589080 513418 589262 513654
rect 589498 513418 589680 513654
rect 589080 513334 589680 513418
rect 589080 513098 589262 513334
rect 589498 513098 589680 513334
rect 589080 477654 589680 513098
rect 589080 477418 589262 477654
rect 589498 477418 589680 477654
rect 589080 477334 589680 477418
rect 589080 477098 589262 477334
rect 589498 477098 589680 477334
rect 589080 441654 589680 477098
rect 589080 441418 589262 441654
rect 589498 441418 589680 441654
rect 589080 441334 589680 441418
rect 589080 441098 589262 441334
rect 589498 441098 589680 441334
rect 589080 405654 589680 441098
rect 589080 405418 589262 405654
rect 589498 405418 589680 405654
rect 589080 405334 589680 405418
rect 589080 405098 589262 405334
rect 589498 405098 589680 405334
rect 589080 369654 589680 405098
rect 589080 369418 589262 369654
rect 589498 369418 589680 369654
rect 589080 369334 589680 369418
rect 589080 369098 589262 369334
rect 589498 369098 589680 369334
rect 589080 333654 589680 369098
rect 589080 333418 589262 333654
rect 589498 333418 589680 333654
rect 589080 333334 589680 333418
rect 589080 333098 589262 333334
rect 589498 333098 589680 333334
rect 589080 297654 589680 333098
rect 589080 297418 589262 297654
rect 589498 297418 589680 297654
rect 589080 297334 589680 297418
rect 589080 297098 589262 297334
rect 589498 297098 589680 297334
rect 589080 261654 589680 297098
rect 589080 261418 589262 261654
rect 589498 261418 589680 261654
rect 589080 261334 589680 261418
rect 589080 261098 589262 261334
rect 589498 261098 589680 261334
rect 589080 225654 589680 261098
rect 589080 225418 589262 225654
rect 589498 225418 589680 225654
rect 589080 225334 589680 225418
rect 589080 225098 589262 225334
rect 589498 225098 589680 225334
rect 589080 189654 589680 225098
rect 589080 189418 589262 189654
rect 589498 189418 589680 189654
rect 589080 189334 589680 189418
rect 589080 189098 589262 189334
rect 589498 189098 589680 189334
rect 589080 153654 589680 189098
rect 589080 153418 589262 153654
rect 589498 153418 589680 153654
rect 589080 153334 589680 153418
rect 589080 153098 589262 153334
rect 589498 153098 589680 153334
rect 589080 117654 589680 153098
rect 589080 117418 589262 117654
rect 589498 117418 589680 117654
rect 589080 117334 589680 117418
rect 589080 117098 589262 117334
rect 589498 117098 589680 117334
rect 589080 81654 589680 117098
rect 589080 81418 589262 81654
rect 589498 81418 589680 81654
rect 589080 81334 589680 81418
rect 589080 81098 589262 81334
rect 589498 81098 589680 81334
rect 589080 45654 589680 81098
rect 589080 45418 589262 45654
rect 589498 45418 589680 45654
rect 589080 45334 589680 45418
rect 589080 45098 589262 45334
rect 589498 45098 589680 45334
rect 589080 9654 589680 45098
rect 589080 9418 589262 9654
rect 589498 9418 589680 9654
rect 589080 9334 589680 9418
rect 589080 9098 589262 9334
rect 589498 9098 589680 9334
rect 589080 -4106 589680 9098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 675654 590620 708982
rect 590020 675418 590202 675654
rect 590438 675418 590620 675654
rect 590020 675334 590620 675418
rect 590020 675098 590202 675334
rect 590438 675098 590620 675334
rect 590020 639654 590620 675098
rect 590020 639418 590202 639654
rect 590438 639418 590620 639654
rect 590020 639334 590620 639418
rect 590020 639098 590202 639334
rect 590438 639098 590620 639334
rect 590020 603654 590620 639098
rect 590020 603418 590202 603654
rect 590438 603418 590620 603654
rect 590020 603334 590620 603418
rect 590020 603098 590202 603334
rect 590438 603098 590620 603334
rect 590020 567654 590620 603098
rect 590020 567418 590202 567654
rect 590438 567418 590620 567654
rect 590020 567334 590620 567418
rect 590020 567098 590202 567334
rect 590438 567098 590620 567334
rect 590020 531654 590620 567098
rect 590020 531418 590202 531654
rect 590438 531418 590620 531654
rect 590020 531334 590620 531418
rect 590020 531098 590202 531334
rect 590438 531098 590620 531334
rect 590020 495654 590620 531098
rect 590020 495418 590202 495654
rect 590438 495418 590620 495654
rect 590020 495334 590620 495418
rect 590020 495098 590202 495334
rect 590438 495098 590620 495334
rect 590020 459654 590620 495098
rect 590020 459418 590202 459654
rect 590438 459418 590620 459654
rect 590020 459334 590620 459418
rect 590020 459098 590202 459334
rect 590438 459098 590620 459334
rect 590020 423654 590620 459098
rect 590020 423418 590202 423654
rect 590438 423418 590620 423654
rect 590020 423334 590620 423418
rect 590020 423098 590202 423334
rect 590438 423098 590620 423334
rect 590020 387654 590620 423098
rect 590020 387418 590202 387654
rect 590438 387418 590620 387654
rect 590020 387334 590620 387418
rect 590020 387098 590202 387334
rect 590438 387098 590620 387334
rect 590020 351654 590620 387098
rect 590020 351418 590202 351654
rect 590438 351418 590620 351654
rect 590020 351334 590620 351418
rect 590020 351098 590202 351334
rect 590438 351098 590620 351334
rect 590020 315654 590620 351098
rect 590020 315418 590202 315654
rect 590438 315418 590620 315654
rect 590020 315334 590620 315418
rect 590020 315098 590202 315334
rect 590438 315098 590620 315334
rect 590020 279654 590620 315098
rect 590020 279418 590202 279654
rect 590438 279418 590620 279654
rect 590020 279334 590620 279418
rect 590020 279098 590202 279334
rect 590438 279098 590620 279334
rect 590020 243654 590620 279098
rect 590020 243418 590202 243654
rect 590438 243418 590620 243654
rect 590020 243334 590620 243418
rect 590020 243098 590202 243334
rect 590438 243098 590620 243334
rect 590020 207654 590620 243098
rect 590020 207418 590202 207654
rect 590438 207418 590620 207654
rect 590020 207334 590620 207418
rect 590020 207098 590202 207334
rect 590438 207098 590620 207334
rect 590020 171654 590620 207098
rect 590020 171418 590202 171654
rect 590438 171418 590620 171654
rect 590020 171334 590620 171418
rect 590020 171098 590202 171334
rect 590438 171098 590620 171334
rect 590020 135654 590620 171098
rect 590020 135418 590202 135654
rect 590438 135418 590620 135654
rect 590020 135334 590620 135418
rect 590020 135098 590202 135334
rect 590438 135098 590620 135334
rect 590020 99654 590620 135098
rect 590020 99418 590202 99654
rect 590438 99418 590620 99654
rect 590020 99334 590620 99418
rect 590020 99098 590202 99334
rect 590438 99098 590620 99334
rect 590020 63654 590620 99098
rect 590020 63418 590202 63654
rect 590438 63418 590620 63654
rect 590020 63334 590620 63418
rect 590020 63098 590202 63334
rect 590438 63098 590620 63334
rect 590020 27654 590620 63098
rect 590020 27418 590202 27654
rect 590438 27418 590620 27654
rect 590020 27334 590620 27418
rect 590020 27098 590202 27334
rect 590438 27098 590620 27334
rect 590020 -5046 590620 27098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 697254 591560 709922
rect 590960 697018 591142 697254
rect 591378 697018 591560 697254
rect 590960 696934 591560 697018
rect 590960 696698 591142 696934
rect 591378 696698 591560 696934
rect 590960 661254 591560 696698
rect 590960 661018 591142 661254
rect 591378 661018 591560 661254
rect 590960 660934 591560 661018
rect 590960 660698 591142 660934
rect 591378 660698 591560 660934
rect 590960 625254 591560 660698
rect 590960 625018 591142 625254
rect 591378 625018 591560 625254
rect 590960 624934 591560 625018
rect 590960 624698 591142 624934
rect 591378 624698 591560 624934
rect 590960 589254 591560 624698
rect 590960 589018 591142 589254
rect 591378 589018 591560 589254
rect 590960 588934 591560 589018
rect 590960 588698 591142 588934
rect 591378 588698 591560 588934
rect 590960 553254 591560 588698
rect 590960 553018 591142 553254
rect 591378 553018 591560 553254
rect 590960 552934 591560 553018
rect 590960 552698 591142 552934
rect 591378 552698 591560 552934
rect 590960 517254 591560 552698
rect 590960 517018 591142 517254
rect 591378 517018 591560 517254
rect 590960 516934 591560 517018
rect 590960 516698 591142 516934
rect 591378 516698 591560 516934
rect 590960 481254 591560 516698
rect 590960 481018 591142 481254
rect 591378 481018 591560 481254
rect 590960 480934 591560 481018
rect 590960 480698 591142 480934
rect 591378 480698 591560 480934
rect 590960 445254 591560 480698
rect 590960 445018 591142 445254
rect 591378 445018 591560 445254
rect 590960 444934 591560 445018
rect 590960 444698 591142 444934
rect 591378 444698 591560 444934
rect 590960 409254 591560 444698
rect 590960 409018 591142 409254
rect 591378 409018 591560 409254
rect 590960 408934 591560 409018
rect 590960 408698 591142 408934
rect 591378 408698 591560 408934
rect 590960 373254 591560 408698
rect 590960 373018 591142 373254
rect 591378 373018 591560 373254
rect 590960 372934 591560 373018
rect 590960 372698 591142 372934
rect 591378 372698 591560 372934
rect 590960 337254 591560 372698
rect 590960 337018 591142 337254
rect 591378 337018 591560 337254
rect 590960 336934 591560 337018
rect 590960 336698 591142 336934
rect 591378 336698 591560 336934
rect 590960 301254 591560 336698
rect 590960 301018 591142 301254
rect 591378 301018 591560 301254
rect 590960 300934 591560 301018
rect 590960 300698 591142 300934
rect 591378 300698 591560 300934
rect 590960 265254 591560 300698
rect 590960 265018 591142 265254
rect 591378 265018 591560 265254
rect 590960 264934 591560 265018
rect 590960 264698 591142 264934
rect 591378 264698 591560 264934
rect 590960 229254 591560 264698
rect 590960 229018 591142 229254
rect 591378 229018 591560 229254
rect 590960 228934 591560 229018
rect 590960 228698 591142 228934
rect 591378 228698 591560 228934
rect 590960 193254 591560 228698
rect 590960 193018 591142 193254
rect 591378 193018 591560 193254
rect 590960 192934 591560 193018
rect 590960 192698 591142 192934
rect 591378 192698 591560 192934
rect 590960 157254 591560 192698
rect 590960 157018 591142 157254
rect 591378 157018 591560 157254
rect 590960 156934 591560 157018
rect 590960 156698 591142 156934
rect 591378 156698 591560 156934
rect 590960 121254 591560 156698
rect 590960 121018 591142 121254
rect 591378 121018 591560 121254
rect 590960 120934 591560 121018
rect 590960 120698 591142 120934
rect 591378 120698 591560 120934
rect 590960 85254 591560 120698
rect 590960 85018 591142 85254
rect 591378 85018 591560 85254
rect 590960 84934 591560 85018
rect 590960 84698 591142 84934
rect 591378 84698 591560 84934
rect 590960 49254 591560 84698
rect 590960 49018 591142 49254
rect 591378 49018 591560 49254
rect 590960 48934 591560 49018
rect 590960 48698 591142 48934
rect 591378 48698 591560 48934
rect 590960 13254 591560 48698
rect 590960 13018 591142 13254
rect 591378 13018 591560 13254
rect 590960 12934 591560 13018
rect 590960 12698 591142 12934
rect 591378 12698 591560 12934
rect 590960 -5986 591560 12698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 679254 592500 710862
rect 591900 679018 592082 679254
rect 592318 679018 592500 679254
rect 591900 678934 592500 679018
rect 591900 678698 592082 678934
rect 592318 678698 592500 678934
rect 591900 643254 592500 678698
rect 591900 643018 592082 643254
rect 592318 643018 592500 643254
rect 591900 642934 592500 643018
rect 591900 642698 592082 642934
rect 592318 642698 592500 642934
rect 591900 607254 592500 642698
rect 591900 607018 592082 607254
rect 592318 607018 592500 607254
rect 591900 606934 592500 607018
rect 591900 606698 592082 606934
rect 592318 606698 592500 606934
rect 591900 571254 592500 606698
rect 591900 571018 592082 571254
rect 592318 571018 592500 571254
rect 591900 570934 592500 571018
rect 591900 570698 592082 570934
rect 592318 570698 592500 570934
rect 591900 535254 592500 570698
rect 591900 535018 592082 535254
rect 592318 535018 592500 535254
rect 591900 534934 592500 535018
rect 591900 534698 592082 534934
rect 592318 534698 592500 534934
rect 591900 499254 592500 534698
rect 591900 499018 592082 499254
rect 592318 499018 592500 499254
rect 591900 498934 592500 499018
rect 591900 498698 592082 498934
rect 592318 498698 592500 498934
rect 591900 463254 592500 498698
rect 591900 463018 592082 463254
rect 592318 463018 592500 463254
rect 591900 462934 592500 463018
rect 591900 462698 592082 462934
rect 592318 462698 592500 462934
rect 591900 427254 592500 462698
rect 591900 427018 592082 427254
rect 592318 427018 592500 427254
rect 591900 426934 592500 427018
rect 591900 426698 592082 426934
rect 592318 426698 592500 426934
rect 591900 391254 592500 426698
rect 591900 391018 592082 391254
rect 592318 391018 592500 391254
rect 591900 390934 592500 391018
rect 591900 390698 592082 390934
rect 592318 390698 592500 390934
rect 591900 355254 592500 390698
rect 591900 355018 592082 355254
rect 592318 355018 592500 355254
rect 591900 354934 592500 355018
rect 591900 354698 592082 354934
rect 592318 354698 592500 354934
rect 591900 319254 592500 354698
rect 591900 319018 592082 319254
rect 592318 319018 592500 319254
rect 591900 318934 592500 319018
rect 591900 318698 592082 318934
rect 592318 318698 592500 318934
rect 591900 283254 592500 318698
rect 591900 283018 592082 283254
rect 592318 283018 592500 283254
rect 591900 282934 592500 283018
rect 591900 282698 592082 282934
rect 592318 282698 592500 282934
rect 591900 247254 592500 282698
rect 591900 247018 592082 247254
rect 592318 247018 592500 247254
rect 591900 246934 592500 247018
rect 591900 246698 592082 246934
rect 592318 246698 592500 246934
rect 591900 211254 592500 246698
rect 591900 211018 592082 211254
rect 592318 211018 592500 211254
rect 591900 210934 592500 211018
rect 591900 210698 592082 210934
rect 592318 210698 592500 210934
rect 591900 175254 592500 210698
rect 591900 175018 592082 175254
rect 592318 175018 592500 175254
rect 591900 174934 592500 175018
rect 591900 174698 592082 174934
rect 592318 174698 592500 174934
rect 591900 139254 592500 174698
rect 591900 139018 592082 139254
rect 592318 139018 592500 139254
rect 591900 138934 592500 139018
rect 591900 138698 592082 138934
rect 592318 138698 592500 138934
rect 591900 103254 592500 138698
rect 591900 103018 592082 103254
rect 592318 103018 592500 103254
rect 591900 102934 592500 103018
rect 591900 102698 592082 102934
rect 592318 102698 592500 102934
rect 591900 67254 592500 102698
rect 591900 67018 592082 67254
rect 592318 67018 592500 67254
rect 591900 66934 592500 67018
rect 591900 66698 592082 66934
rect 592318 66698 592500 66934
rect 591900 31254 592500 66698
rect 591900 31018 592082 31254
rect 592318 31018 592500 31254
rect 591900 30934 592500 31018
rect 591900 30698 592082 30934
rect 592318 30698 592500 30934
rect 569604 -7162 569786 -6926
rect 570022 -7162 570204 -6926
rect 569604 -7246 570204 -7162
rect 569604 -7482 569786 -7246
rect 570022 -7482 570204 -7246
rect 569604 -7504 570204 -7482
rect 591900 -6926 592500 30698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 679018 -8158 679254
rect -8394 678698 -8158 678934
rect -8394 643018 -8158 643254
rect -8394 642698 -8158 642934
rect -8394 607018 -8158 607254
rect -8394 606698 -8158 606934
rect -8394 571018 -8158 571254
rect -8394 570698 -8158 570934
rect -8394 535018 -8158 535254
rect -8394 534698 -8158 534934
rect -8394 499018 -8158 499254
rect -8394 498698 -8158 498934
rect -8394 463018 -8158 463254
rect -8394 462698 -8158 462934
rect -8394 427018 -8158 427254
rect -8394 426698 -8158 426934
rect -8394 391018 -8158 391254
rect -8394 390698 -8158 390934
rect -8394 355018 -8158 355254
rect -8394 354698 -8158 354934
rect -8394 319018 -8158 319254
rect -8394 318698 -8158 318934
rect -8394 283018 -8158 283254
rect -8394 282698 -8158 282934
rect -8394 247018 -8158 247254
rect -8394 246698 -8158 246934
rect -8394 211018 -8158 211254
rect -8394 210698 -8158 210934
rect -8394 175018 -8158 175254
rect -8394 174698 -8158 174934
rect -8394 139018 -8158 139254
rect -8394 138698 -8158 138934
rect -8394 103018 -8158 103254
rect -8394 102698 -8158 102934
rect -8394 67018 -8158 67254
rect -8394 66698 -8158 66934
rect -8394 31018 -8158 31254
rect -8394 30698 -8158 30934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 11786 710242 12022 710478
rect 11786 709922 12022 710158
rect -7454 697018 -7218 697254
rect -7454 696698 -7218 696934
rect -7454 661018 -7218 661254
rect -7454 660698 -7218 660934
rect -7454 625018 -7218 625254
rect -7454 624698 -7218 624934
rect -7454 589018 -7218 589254
rect -7454 588698 -7218 588934
rect -7454 553018 -7218 553254
rect -7454 552698 -7218 552934
rect -7454 517018 -7218 517254
rect -7454 516698 -7218 516934
rect -7454 481018 -7218 481254
rect -7454 480698 -7218 480934
rect -7454 445018 -7218 445254
rect -7454 444698 -7218 444934
rect -7454 409018 -7218 409254
rect -7454 408698 -7218 408934
rect -7454 373018 -7218 373254
rect -7454 372698 -7218 372934
rect -7454 337018 -7218 337254
rect -7454 336698 -7218 336934
rect -7454 301018 -7218 301254
rect -7454 300698 -7218 300934
rect -7454 265018 -7218 265254
rect -7454 264698 -7218 264934
rect -7454 229018 -7218 229254
rect -7454 228698 -7218 228934
rect -7454 193018 -7218 193254
rect -7454 192698 -7218 192934
rect -7454 157018 -7218 157254
rect -7454 156698 -7218 156934
rect -7454 121018 -7218 121254
rect -7454 120698 -7218 120934
rect -7454 85018 -7218 85254
rect -7454 84698 -7218 84934
rect -7454 49018 -7218 49254
rect -7454 48698 -7218 48934
rect -7454 13018 -7218 13254
rect -7454 12698 -7218 12934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 675418 -6278 675654
rect -6514 675098 -6278 675334
rect -6514 639418 -6278 639654
rect -6514 639098 -6278 639334
rect -6514 603418 -6278 603654
rect -6514 603098 -6278 603334
rect -6514 567418 -6278 567654
rect -6514 567098 -6278 567334
rect -6514 531418 -6278 531654
rect -6514 531098 -6278 531334
rect -6514 495418 -6278 495654
rect -6514 495098 -6278 495334
rect -6514 459418 -6278 459654
rect -6514 459098 -6278 459334
rect -6514 423418 -6278 423654
rect -6514 423098 -6278 423334
rect -6514 387418 -6278 387654
rect -6514 387098 -6278 387334
rect -6514 351418 -6278 351654
rect -6514 351098 -6278 351334
rect -6514 315418 -6278 315654
rect -6514 315098 -6278 315334
rect -6514 279418 -6278 279654
rect -6514 279098 -6278 279334
rect -6514 243418 -6278 243654
rect -6514 243098 -6278 243334
rect -6514 207418 -6278 207654
rect -6514 207098 -6278 207334
rect -6514 171418 -6278 171654
rect -6514 171098 -6278 171334
rect -6514 135418 -6278 135654
rect -6514 135098 -6278 135334
rect -6514 99418 -6278 99654
rect -6514 99098 -6278 99334
rect -6514 63418 -6278 63654
rect -6514 63098 -6278 63334
rect -6514 27418 -6278 27654
rect -6514 27098 -6278 27334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 8186 708362 8422 708598
rect 8186 708042 8422 708278
rect -5574 693418 -5338 693654
rect -5574 693098 -5338 693334
rect -5574 657418 -5338 657654
rect -5574 657098 -5338 657334
rect -5574 621418 -5338 621654
rect -5574 621098 -5338 621334
rect -5574 585418 -5338 585654
rect -5574 585098 -5338 585334
rect -5574 549418 -5338 549654
rect -5574 549098 -5338 549334
rect -5574 513418 -5338 513654
rect -5574 513098 -5338 513334
rect -5574 477418 -5338 477654
rect -5574 477098 -5338 477334
rect -5574 441418 -5338 441654
rect -5574 441098 -5338 441334
rect -5574 405418 -5338 405654
rect -5574 405098 -5338 405334
rect -5574 369418 -5338 369654
rect -5574 369098 -5338 369334
rect -5574 333418 -5338 333654
rect -5574 333098 -5338 333334
rect -5574 297418 -5338 297654
rect -5574 297098 -5338 297334
rect -5574 261418 -5338 261654
rect -5574 261098 -5338 261334
rect -5574 225418 -5338 225654
rect -5574 225098 -5338 225334
rect -5574 189418 -5338 189654
rect -5574 189098 -5338 189334
rect -5574 153418 -5338 153654
rect -5574 153098 -5338 153334
rect -5574 117418 -5338 117654
rect -5574 117098 -5338 117334
rect -5574 81418 -5338 81654
rect -5574 81098 -5338 81334
rect -5574 45418 -5338 45654
rect -5574 45098 -5338 45334
rect -5574 9418 -5338 9654
rect -5574 9098 -5338 9334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 671818 -4398 672054
rect -4634 671498 -4398 671734
rect -4634 635818 -4398 636054
rect -4634 635498 -4398 635734
rect -4634 599818 -4398 600054
rect -4634 599498 -4398 599734
rect -4634 563818 -4398 564054
rect -4634 563498 -4398 563734
rect -4634 527818 -4398 528054
rect -4634 527498 -4398 527734
rect -4634 491818 -4398 492054
rect -4634 491498 -4398 491734
rect -4634 455818 -4398 456054
rect -4634 455498 -4398 455734
rect -4634 419818 -4398 420054
rect -4634 419498 -4398 419734
rect -4634 383818 -4398 384054
rect -4634 383498 -4398 383734
rect -4634 347818 -4398 348054
rect -4634 347498 -4398 347734
rect -4634 311818 -4398 312054
rect -4634 311498 -4398 311734
rect -4634 275818 -4398 276054
rect -4634 275498 -4398 275734
rect -4634 239818 -4398 240054
rect -4634 239498 -4398 239734
rect -4634 203818 -4398 204054
rect -4634 203498 -4398 203734
rect -4634 167818 -4398 168054
rect -4634 167498 -4398 167734
rect -4634 131818 -4398 132054
rect -4634 131498 -4398 131734
rect -4634 95818 -4398 96054
rect -4634 95498 -4398 95734
rect -4634 59818 -4398 60054
rect -4634 59498 -4398 59734
rect -4634 23818 -4398 24054
rect -4634 23498 -4398 23734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 4586 706482 4822 706718
rect 4586 706162 4822 706398
rect -3694 689818 -3458 690054
rect -3694 689498 -3458 689734
rect -3694 653818 -3458 654054
rect -3694 653498 -3458 653734
rect -3694 617818 -3458 618054
rect -3694 617498 -3458 617734
rect -3694 581818 -3458 582054
rect -3694 581498 -3458 581734
rect -3694 545818 -3458 546054
rect -3694 545498 -3458 545734
rect -3694 509818 -3458 510054
rect -3694 509498 -3458 509734
rect -3694 473818 -3458 474054
rect -3694 473498 -3458 473734
rect -3694 437818 -3458 438054
rect -3694 437498 -3458 437734
rect -3694 401818 -3458 402054
rect -3694 401498 -3458 401734
rect -3694 365818 -3458 366054
rect -3694 365498 -3458 365734
rect -3694 329818 -3458 330054
rect -3694 329498 -3458 329734
rect -3694 293818 -3458 294054
rect -3694 293498 -3458 293734
rect -3694 257818 -3458 258054
rect -3694 257498 -3458 257734
rect -3694 221818 -3458 222054
rect -3694 221498 -3458 221734
rect -3694 185818 -3458 186054
rect -3694 185498 -3458 185734
rect -3694 149818 -3458 150054
rect -3694 149498 -3458 149734
rect -3694 113818 -3458 114054
rect -3694 113498 -3458 113734
rect -3694 77818 -3458 78054
rect -3694 77498 -3458 77734
rect -3694 41818 -3458 42054
rect -3694 41498 -3458 41734
rect -3694 5818 -3458 6054
rect -3694 5498 -3458 5734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 4586 -2462 4822 -2226
rect 4586 -2782 4822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 8186 -4342 8422 -4106
rect 8186 -4662 8422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 29786 711182 30022 711418
rect 29786 710862 30022 711098
rect 26186 709302 26422 709538
rect 26186 708982 26422 709218
rect 22586 707422 22822 707658
rect 22586 707102 22822 707338
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3402 22822 -3166
rect 22586 -3722 22822 -3486
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5282 26422 -5046
rect 26186 -5602 26422 -5366
rect 47786 710242 48022 710478
rect 47786 709922 48022 710158
rect 44186 708362 44422 708598
rect 44186 708042 44422 708278
rect 40586 706482 40822 706718
rect 40586 706162 40822 706398
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6222 12022 -5986
rect 11786 -6542 12022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2462 40822 -2226
rect 40586 -2782 40822 -2546
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4342 44422 -4106
rect 44186 -4662 44422 -4426
rect 65786 711182 66022 711418
rect 65786 710862 66022 711098
rect 62186 709302 62422 709538
rect 62186 708982 62422 709218
rect 58586 707422 58822 707658
rect 58586 707102 58822 707338
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7162 30022 -6926
rect 29786 -7482 30022 -7246
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3402 58822 -3166
rect 58586 -3722 58822 -3486
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5282 62422 -5046
rect 62186 -5602 62422 -5366
rect 83786 710242 84022 710478
rect 83786 709922 84022 710158
rect 80186 708362 80422 708598
rect 80186 708042 80422 708278
rect 76586 706482 76822 706718
rect 76586 706162 76822 706398
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6222 48022 -5986
rect 47786 -6542 48022 -6306
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2462 76822 -2226
rect 76586 -2782 76822 -2546
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4342 80422 -4106
rect 80186 -4662 80422 -4426
rect 101786 711182 102022 711418
rect 101786 710862 102022 711098
rect 98186 709302 98422 709538
rect 98186 708982 98422 709218
rect 94586 707422 94822 707658
rect 94586 707102 94822 707338
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 83786 373018 84022 373254
rect 83786 372698 84022 372934
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7162 66022 -6926
rect 65786 -7482 66022 -7246
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3402 94822 -3166
rect 94586 -3722 94822 -3486
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 98186 531418 98422 531654
rect 98186 531098 98422 531334
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 98186 387418 98422 387654
rect 98186 387098 98422 387334
rect 98186 351418 98422 351654
rect 98186 351098 98422 351334
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5282 98422 -5046
rect 98186 -5602 98422 -5366
rect 119786 710242 120022 710478
rect 119786 709922 120022 710158
rect 116186 708362 116422 708598
rect 116186 708042 116422 708278
rect 112586 706482 112822 706718
rect 112586 706162 112822 706398
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 101786 535018 102022 535254
rect 101786 534698 102022 534934
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 101786 391018 102022 391254
rect 101786 390698 102022 390934
rect 101786 355018 102022 355254
rect 101786 354698 102022 354934
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6222 84022 -5986
rect 83786 -6542 84022 -6306
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2462 112822 -2226
rect 112586 -2782 112822 -2546
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 116186 369418 116422 369654
rect 116186 369098 116422 369334
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4342 116422 -4106
rect 116186 -4662 116422 -4426
rect 137786 711182 138022 711418
rect 137786 710862 138022 711098
rect 134186 709302 134422 709538
rect 134186 708982 134422 709218
rect 130586 707422 130822 707658
rect 130586 707102 130822 707338
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 119786 373018 120022 373254
rect 119786 372698 120022 372934
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7162 102022 -6926
rect 101786 -7482 102022 -7246
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3402 130822 -3166
rect 130586 -3722 130822 -3486
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5282 134422 -5046
rect 134186 -5602 134422 -5366
rect 155786 710242 156022 710478
rect 155786 709922 156022 710158
rect 152186 708362 152422 708598
rect 152186 708042 152422 708278
rect 148586 706482 148822 706718
rect 148586 706162 148822 706398
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6222 120022 -5986
rect 119786 -6542 120022 -6306
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2462 148822 -2226
rect 148586 -2782 148822 -2546
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 173786 711182 174022 711418
rect 173786 710862 174022 711098
rect 170186 709302 170422 709538
rect 170186 708982 170422 709218
rect 166586 707422 166822 707658
rect 166586 707102 166822 707338
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 191786 710242 192022 710478
rect 191786 709922 192022 710158
rect 188186 708362 188422 708598
rect 188186 708042 188422 708278
rect 184586 706482 184822 706718
rect 184586 706162 184822 706398
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 209786 711182 210022 711418
rect 209786 710862 210022 711098
rect 206186 709302 206422 709538
rect 206186 708982 206422 709218
rect 202586 707422 202822 707658
rect 202586 707102 202822 707338
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 206186 531418 206422 531654
rect 206186 531098 206422 531334
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 227786 710242 228022 710478
rect 227786 709922 228022 710158
rect 224186 708362 224422 708598
rect 224186 708042 224422 708278
rect 220586 706482 220822 706718
rect 220586 706162 220822 706398
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 209786 535018 210022 535254
rect 209786 534698 210022 534934
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 245786 711182 246022 711418
rect 245786 710862 246022 711098
rect 242186 709302 242422 709538
rect 242186 708982 242422 709218
rect 238586 707422 238822 707658
rect 238586 707102 238822 707338
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 238586 419818 238822 420054
rect 238586 419498 238822 419734
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 242186 423418 242422 423654
rect 242186 423098 242422 423334
rect 263786 710242 264022 710478
rect 263786 709922 264022 710158
rect 260186 708362 260422 708598
rect 260186 708042 260422 708278
rect 256586 706482 256822 706718
rect 256586 706162 256822 706398
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 260186 477418 260422 477654
rect 260186 477098 260422 477334
rect 260186 441418 260422 441654
rect 260186 441098 260422 441334
rect 281786 711182 282022 711418
rect 281786 710862 282022 711098
rect 278186 709302 278422 709538
rect 278186 708982 278422 709218
rect 274586 707422 274822 707658
rect 274586 707102 274822 707338
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 263786 481018 264022 481254
rect 263786 480698 264022 480934
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 274586 419818 274822 420054
rect 274586 419498 274822 419734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 278186 459418 278422 459654
rect 278186 459098 278422 459334
rect 278186 423418 278422 423654
rect 278186 423098 278422 423334
rect 299786 710242 300022 710478
rect 299786 709922 300022 710158
rect 296186 708362 296422 708598
rect 296186 708042 296422 708278
rect 292586 706482 292822 706718
rect 292586 706162 292822 706398
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 281786 463018 282022 463254
rect 281786 462698 282022 462934
rect 281786 427018 282022 427254
rect 281786 426698 282022 426934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 317786 711182 318022 711418
rect 317786 710862 318022 711098
rect 314186 709302 314422 709538
rect 314186 708982 314422 709218
rect 310586 707422 310822 707658
rect 310586 707102 310822 707338
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 314186 567418 314422 567654
rect 314186 567098 314422 567334
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 335786 710242 336022 710478
rect 335786 709922 336022 710158
rect 332186 708362 332422 708598
rect 332186 708042 332422 708278
rect 328586 706482 328822 706718
rect 328586 706162 328822 706398
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 317786 571018 318022 571254
rect 317786 570698 318022 570934
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 353786 711182 354022 711418
rect 353786 710862 354022 711098
rect 350186 709302 350422 709538
rect 350186 708982 350422 709218
rect 346586 707422 346822 707658
rect 346586 707102 346822 707338
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 335786 517018 336022 517254
rect 335786 516698 336022 516934
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 350186 567418 350422 567654
rect 350186 567098 350422 567334
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 371786 710242 372022 710478
rect 371786 709922 372022 710158
rect 368186 708362 368422 708598
rect 368186 708042 368422 708278
rect 364586 706482 364822 706718
rect 364586 706162 364822 706398
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 353786 571018 354022 571254
rect 353786 570698 354022 570934
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 389786 711182 390022 711418
rect 389786 710862 390022 711098
rect 386186 709302 386422 709538
rect 386186 708982 386422 709218
rect 382586 707422 382822 707658
rect 382586 707102 382822 707338
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 371786 517018 372022 517254
rect 371786 516698 372022 516934
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 407786 710242 408022 710478
rect 407786 709922 408022 710158
rect 404186 708362 404422 708598
rect 404186 708042 404422 708278
rect 400586 706482 400822 706718
rect 400586 706162 400822 706398
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4342 152422 -4106
rect 152186 -4662 152422 -4426
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7162 138022 -6926
rect 137786 -7482 138022 -7246
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3402 166822 -3166
rect 166586 -3722 166822 -3486
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5282 170422 -5046
rect 170186 -5602 170422 -5366
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6222 156022 -5986
rect 155786 -6542 156022 -6306
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2462 184822 -2226
rect 184586 -2782 184822 -2546
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4342 188422 -4106
rect 188186 -4662 188422 -4426
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7162 174022 -6926
rect 173786 -7482 174022 -7246
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3402 202822 -3166
rect 202586 -3722 202822 -3486
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5282 206422 -5046
rect 206186 -5602 206422 -5366
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6222 192022 -5986
rect 191786 -6542 192022 -6306
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2462 220822 -2226
rect 220586 -2782 220822 -2546
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4342 224422 -4106
rect 224186 -4662 224422 -4426
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7162 210022 -6926
rect 209786 -7482 210022 -7246
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3402 238822 -3166
rect 238586 -3722 238822 -3486
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5282 242422 -5046
rect 242186 -5602 242422 -5366
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6222 228022 -5986
rect 227786 -6542 228022 -6306
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2462 256822 -2226
rect 256586 -2782 256822 -2546
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4342 260422 -4106
rect 260186 -4662 260422 -4426
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7162 246022 -6926
rect 245786 -7482 246022 -7246
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3402 274822 -3166
rect 274586 -3722 274822 -3486
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5282 278422 -5046
rect 278186 -5602 278422 -5366
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6222 264022 -5986
rect 263786 -6542 264022 -6306
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2462 292822 -2226
rect 292586 -2782 292822 -2546
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4342 296422 -4106
rect 296186 -4662 296422 -4426
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7162 282022 -6926
rect 281786 -7482 282022 -7246
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3402 310822 -3166
rect 310586 -3722 310822 -3486
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5282 314422 -5046
rect 314186 -5602 314422 -5366
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6222 300022 -5986
rect 299786 -6542 300022 -6306
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2462 328822 -2226
rect 328586 -2782 328822 -2546
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4342 332422 -4106
rect 332186 -4662 332422 -4426
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7162 318022 -6926
rect 317786 -7482 318022 -7246
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3402 346822 -3166
rect 346586 -3722 346822 -3486
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5282 350422 -5046
rect 350186 -5602 350422 -5366
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6222 336022 -5986
rect 335786 -6542 336022 -6306
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2462 364822 -2226
rect 364586 -2782 364822 -2546
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4342 368422 -4106
rect 368186 -4662 368422 -4426
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7162 354022 -6926
rect 353786 -7482 354022 -7246
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3402 382822 -3166
rect 382586 -3722 382822 -3486
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5282 386422 -5046
rect 386186 -5602 386422 -5366
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6222 372022 -5986
rect 371786 -6542 372022 -6306
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 400586 365818 400822 366054
rect 400586 365498 400822 365734
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2462 400822 -2226
rect 400586 -2782 400822 -2546
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 404186 369418 404422 369654
rect 404186 369098 404422 369334
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4342 404422 -4106
rect 404186 -4662 404422 -4426
rect 425786 711182 426022 711418
rect 425786 710862 426022 711098
rect 422186 709302 422422 709538
rect 422186 708982 422422 709218
rect 418586 707422 418822 707658
rect 418586 707102 418822 707338
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 407786 373018 408022 373254
rect 407786 372698 408022 372934
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7162 390022 -6926
rect 389786 -7482 390022 -7246
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3402 418822 -3166
rect 418586 -3722 418822 -3486
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5282 422422 -5046
rect 422186 -5602 422422 -5366
rect 443786 710242 444022 710478
rect 443786 709922 444022 710158
rect 440186 708362 440422 708598
rect 440186 708042 440422 708278
rect 436586 706482 436822 706718
rect 436586 706162 436822 706398
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6222 408022 -5986
rect 407786 -6542 408022 -6306
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2462 436822 -2226
rect 436586 -2782 436822 -2546
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4342 440422 -4106
rect 440186 -4662 440422 -4426
rect 461786 711182 462022 711418
rect 461786 710862 462022 711098
rect 458186 709302 458422 709538
rect 458186 708982 458422 709218
rect 454586 707422 454822 707658
rect 454586 707102 454822 707338
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7162 426022 -6926
rect 425786 -7482 426022 -7246
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3402 454822 -3166
rect 454586 -3722 454822 -3486
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5282 458422 -5046
rect 458186 -5602 458422 -5366
rect 479786 710242 480022 710478
rect 479786 709922 480022 710158
rect 476186 708362 476422 708598
rect 476186 708042 476422 708278
rect 472586 706482 472822 706718
rect 472586 706162 472822 706398
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6222 444022 -5986
rect 443786 -6542 444022 -6306
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2462 472822 -2226
rect 472586 -2782 472822 -2546
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4342 476422 -4106
rect 476186 -4662 476422 -4426
rect 497786 711182 498022 711418
rect 497786 710862 498022 711098
rect 494186 709302 494422 709538
rect 494186 708982 494422 709218
rect 490586 707422 490822 707658
rect 490586 707102 490822 707338
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7162 462022 -6926
rect 461786 -7482 462022 -7246
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3402 490822 -3166
rect 490586 -3722 490822 -3486
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5282 494422 -5046
rect 494186 -5602 494422 -5366
rect 515786 710242 516022 710478
rect 515786 709922 516022 710158
rect 512186 708362 512422 708598
rect 512186 708042 512422 708278
rect 508586 706482 508822 706718
rect 508586 706162 508822 706398
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6222 480022 -5986
rect 479786 -6542 480022 -6306
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2462 508822 -2226
rect 508586 -2782 508822 -2546
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4342 512422 -4106
rect 512186 -4662 512422 -4426
rect 533786 711182 534022 711418
rect 533786 710862 534022 711098
rect 530186 709302 530422 709538
rect 530186 708982 530422 709218
rect 526586 707422 526822 707658
rect 526586 707102 526822 707338
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7162 498022 -6926
rect 497786 -7482 498022 -7246
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3402 526822 -3166
rect 526586 -3722 526822 -3486
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5282 530422 -5046
rect 530186 -5602 530422 -5366
rect 551786 710242 552022 710478
rect 551786 709922 552022 710158
rect 548186 708362 548422 708598
rect 548186 708042 548422 708278
rect 544586 706482 544822 706718
rect 544586 706162 544822 706398
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6222 516022 -5986
rect 515786 -6542 516022 -6306
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2462 544822 -2226
rect 544586 -2782 544822 -2546
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4342 548422 -4106
rect 548186 -4662 548422 -4426
rect 569786 711182 570022 711418
rect 569786 710862 570022 711098
rect 566186 709302 566422 709538
rect 566186 708982 566422 709218
rect 562586 707422 562822 707658
rect 562586 707102 562822 707338
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7162 534022 -6926
rect 533786 -7482 534022 -7246
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3402 562822 -3166
rect 562586 -3722 562822 -3486
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5282 566422 -5046
rect 566186 -5602 566422 -5366
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 580586 706482 580822 706718
rect 580586 706162 580822 706398
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6222 552022 -5986
rect 551786 -6542 552022 -6306
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 689818 587618 690054
rect 587382 689498 587618 689734
rect 587382 653818 587618 654054
rect 587382 653498 587618 653734
rect 587382 617818 587618 618054
rect 587382 617498 587618 617734
rect 587382 581818 587618 582054
rect 587382 581498 587618 581734
rect 587382 545818 587618 546054
rect 587382 545498 587618 545734
rect 587382 509818 587618 510054
rect 587382 509498 587618 509734
rect 587382 473818 587618 474054
rect 587382 473498 587618 473734
rect 587382 437818 587618 438054
rect 587382 437498 587618 437734
rect 587382 401818 587618 402054
rect 587382 401498 587618 401734
rect 587382 365818 587618 366054
rect 587382 365498 587618 365734
rect 587382 329818 587618 330054
rect 587382 329498 587618 329734
rect 587382 293818 587618 294054
rect 587382 293498 587618 293734
rect 587382 257818 587618 258054
rect 587382 257498 587618 257734
rect 587382 221818 587618 222054
rect 587382 221498 587618 221734
rect 587382 185818 587618 186054
rect 587382 185498 587618 185734
rect 587382 149818 587618 150054
rect 587382 149498 587618 149734
rect 587382 113818 587618 114054
rect 587382 113498 587618 113734
rect 587382 77818 587618 78054
rect 587382 77498 587618 77734
rect 587382 41818 587618 42054
rect 587382 41498 587618 41734
rect 587382 5818 587618 6054
rect 587382 5498 587618 5734
rect 580586 -2462 580822 -2226
rect 580586 -2782 580822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 671818 588558 672054
rect 588322 671498 588558 671734
rect 588322 635818 588558 636054
rect 588322 635498 588558 635734
rect 588322 599818 588558 600054
rect 588322 599498 588558 599734
rect 588322 563818 588558 564054
rect 588322 563498 588558 563734
rect 588322 527818 588558 528054
rect 588322 527498 588558 527734
rect 588322 491818 588558 492054
rect 588322 491498 588558 491734
rect 588322 455818 588558 456054
rect 588322 455498 588558 455734
rect 588322 419818 588558 420054
rect 588322 419498 588558 419734
rect 588322 383818 588558 384054
rect 588322 383498 588558 383734
rect 588322 347818 588558 348054
rect 588322 347498 588558 347734
rect 588322 311818 588558 312054
rect 588322 311498 588558 311734
rect 588322 275818 588558 276054
rect 588322 275498 588558 275734
rect 588322 239818 588558 240054
rect 588322 239498 588558 239734
rect 588322 203818 588558 204054
rect 588322 203498 588558 203734
rect 588322 167818 588558 168054
rect 588322 167498 588558 167734
rect 588322 131818 588558 132054
rect 588322 131498 588558 131734
rect 588322 95818 588558 96054
rect 588322 95498 588558 95734
rect 588322 59818 588558 60054
rect 588322 59498 588558 59734
rect 588322 23818 588558 24054
rect 588322 23498 588558 23734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 693418 589498 693654
rect 589262 693098 589498 693334
rect 589262 657418 589498 657654
rect 589262 657098 589498 657334
rect 589262 621418 589498 621654
rect 589262 621098 589498 621334
rect 589262 585418 589498 585654
rect 589262 585098 589498 585334
rect 589262 549418 589498 549654
rect 589262 549098 589498 549334
rect 589262 513418 589498 513654
rect 589262 513098 589498 513334
rect 589262 477418 589498 477654
rect 589262 477098 589498 477334
rect 589262 441418 589498 441654
rect 589262 441098 589498 441334
rect 589262 405418 589498 405654
rect 589262 405098 589498 405334
rect 589262 369418 589498 369654
rect 589262 369098 589498 369334
rect 589262 333418 589498 333654
rect 589262 333098 589498 333334
rect 589262 297418 589498 297654
rect 589262 297098 589498 297334
rect 589262 261418 589498 261654
rect 589262 261098 589498 261334
rect 589262 225418 589498 225654
rect 589262 225098 589498 225334
rect 589262 189418 589498 189654
rect 589262 189098 589498 189334
rect 589262 153418 589498 153654
rect 589262 153098 589498 153334
rect 589262 117418 589498 117654
rect 589262 117098 589498 117334
rect 589262 81418 589498 81654
rect 589262 81098 589498 81334
rect 589262 45418 589498 45654
rect 589262 45098 589498 45334
rect 589262 9418 589498 9654
rect 589262 9098 589498 9334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 675418 590438 675654
rect 590202 675098 590438 675334
rect 590202 639418 590438 639654
rect 590202 639098 590438 639334
rect 590202 603418 590438 603654
rect 590202 603098 590438 603334
rect 590202 567418 590438 567654
rect 590202 567098 590438 567334
rect 590202 531418 590438 531654
rect 590202 531098 590438 531334
rect 590202 495418 590438 495654
rect 590202 495098 590438 495334
rect 590202 459418 590438 459654
rect 590202 459098 590438 459334
rect 590202 423418 590438 423654
rect 590202 423098 590438 423334
rect 590202 387418 590438 387654
rect 590202 387098 590438 387334
rect 590202 351418 590438 351654
rect 590202 351098 590438 351334
rect 590202 315418 590438 315654
rect 590202 315098 590438 315334
rect 590202 279418 590438 279654
rect 590202 279098 590438 279334
rect 590202 243418 590438 243654
rect 590202 243098 590438 243334
rect 590202 207418 590438 207654
rect 590202 207098 590438 207334
rect 590202 171418 590438 171654
rect 590202 171098 590438 171334
rect 590202 135418 590438 135654
rect 590202 135098 590438 135334
rect 590202 99418 590438 99654
rect 590202 99098 590438 99334
rect 590202 63418 590438 63654
rect 590202 63098 590438 63334
rect 590202 27418 590438 27654
rect 590202 27098 590438 27334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 697018 591378 697254
rect 591142 696698 591378 696934
rect 591142 661018 591378 661254
rect 591142 660698 591378 660934
rect 591142 625018 591378 625254
rect 591142 624698 591378 624934
rect 591142 589018 591378 589254
rect 591142 588698 591378 588934
rect 591142 553018 591378 553254
rect 591142 552698 591378 552934
rect 591142 517018 591378 517254
rect 591142 516698 591378 516934
rect 591142 481018 591378 481254
rect 591142 480698 591378 480934
rect 591142 445018 591378 445254
rect 591142 444698 591378 444934
rect 591142 409018 591378 409254
rect 591142 408698 591378 408934
rect 591142 373018 591378 373254
rect 591142 372698 591378 372934
rect 591142 337018 591378 337254
rect 591142 336698 591378 336934
rect 591142 301018 591378 301254
rect 591142 300698 591378 300934
rect 591142 265018 591378 265254
rect 591142 264698 591378 264934
rect 591142 229018 591378 229254
rect 591142 228698 591378 228934
rect 591142 193018 591378 193254
rect 591142 192698 591378 192934
rect 591142 157018 591378 157254
rect 591142 156698 591378 156934
rect 591142 121018 591378 121254
rect 591142 120698 591378 120934
rect 591142 85018 591378 85254
rect 591142 84698 591378 84934
rect 591142 49018 591378 49254
rect 591142 48698 591378 48934
rect 591142 13018 591378 13254
rect 591142 12698 591378 12934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 679018 592318 679254
rect 592082 678698 592318 678934
rect 592082 643018 592318 643254
rect 592082 642698 592318 642934
rect 592082 607018 592318 607254
rect 592082 606698 592318 606934
rect 592082 571018 592318 571254
rect 592082 570698 592318 570934
rect 592082 535018 592318 535254
rect 592082 534698 592318 534934
rect 592082 499018 592318 499254
rect 592082 498698 592318 498934
rect 592082 463018 592318 463254
rect 592082 462698 592318 462934
rect 592082 427018 592318 427254
rect 592082 426698 592318 426934
rect 592082 391018 592318 391254
rect 592082 390698 592318 390934
rect 592082 355018 592318 355254
rect 592082 354698 592318 354934
rect 592082 319018 592318 319254
rect 592082 318698 592318 318934
rect 592082 283018 592318 283254
rect 592082 282698 592318 282934
rect 592082 247018 592318 247254
rect 592082 246698 592318 246934
rect 592082 211018 592318 211254
rect 592082 210698 592318 210934
rect 592082 175018 592318 175254
rect 592082 174698 592318 174934
rect 592082 139018 592318 139254
rect 592082 138698 592318 138934
rect 592082 103018 592318 103254
rect 592082 102698 592318 102934
rect 592082 67018 592318 67254
rect 592082 66698 592318 66934
rect 592082 31018 592318 31254
rect 592082 30698 592318 30934
rect 569786 -7162 570022 -6926
rect 569786 -7482 570022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 29786 711418
rect 30022 711182 65786 711418
rect 66022 711182 101786 711418
rect 102022 711182 137786 711418
rect 138022 711182 173786 711418
rect 174022 711182 209786 711418
rect 210022 711182 245786 711418
rect 246022 711182 281786 711418
rect 282022 711182 317786 711418
rect 318022 711182 353786 711418
rect 354022 711182 389786 711418
rect 390022 711182 425786 711418
rect 426022 711182 461786 711418
rect 462022 711182 497786 711418
rect 498022 711182 533786 711418
rect 534022 711182 569786 711418
rect 570022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 29786 711098
rect 30022 710862 65786 711098
rect 66022 710862 101786 711098
rect 102022 710862 137786 711098
rect 138022 710862 173786 711098
rect 174022 710862 209786 711098
rect 210022 710862 245786 711098
rect 246022 710862 281786 711098
rect 282022 710862 317786 711098
rect 318022 710862 353786 711098
rect 354022 710862 389786 711098
rect 390022 710862 425786 711098
rect 426022 710862 461786 711098
rect 462022 710862 497786 711098
rect 498022 710862 533786 711098
rect 534022 710862 569786 711098
rect 570022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 11786 710478
rect 12022 710242 47786 710478
rect 48022 710242 83786 710478
rect 84022 710242 119786 710478
rect 120022 710242 155786 710478
rect 156022 710242 191786 710478
rect 192022 710242 227786 710478
rect 228022 710242 263786 710478
rect 264022 710242 299786 710478
rect 300022 710242 335786 710478
rect 336022 710242 371786 710478
rect 372022 710242 407786 710478
rect 408022 710242 443786 710478
rect 444022 710242 479786 710478
rect 480022 710242 515786 710478
rect 516022 710242 551786 710478
rect 552022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 11786 710158
rect 12022 709922 47786 710158
rect 48022 709922 83786 710158
rect 84022 709922 119786 710158
rect 120022 709922 155786 710158
rect 156022 709922 191786 710158
rect 192022 709922 227786 710158
rect 228022 709922 263786 710158
rect 264022 709922 299786 710158
rect 300022 709922 335786 710158
rect 336022 709922 371786 710158
rect 372022 709922 407786 710158
rect 408022 709922 443786 710158
rect 444022 709922 479786 710158
rect 480022 709922 515786 710158
rect 516022 709922 551786 710158
rect 552022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 26186 709538
rect 26422 709302 62186 709538
rect 62422 709302 98186 709538
rect 98422 709302 134186 709538
rect 134422 709302 170186 709538
rect 170422 709302 206186 709538
rect 206422 709302 242186 709538
rect 242422 709302 278186 709538
rect 278422 709302 314186 709538
rect 314422 709302 350186 709538
rect 350422 709302 386186 709538
rect 386422 709302 422186 709538
rect 422422 709302 458186 709538
rect 458422 709302 494186 709538
rect 494422 709302 530186 709538
rect 530422 709302 566186 709538
rect 566422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 26186 709218
rect 26422 708982 62186 709218
rect 62422 708982 98186 709218
rect 98422 708982 134186 709218
rect 134422 708982 170186 709218
rect 170422 708982 206186 709218
rect 206422 708982 242186 709218
rect 242422 708982 278186 709218
rect 278422 708982 314186 709218
rect 314422 708982 350186 709218
rect 350422 708982 386186 709218
rect 386422 708982 422186 709218
rect 422422 708982 458186 709218
rect 458422 708982 494186 709218
rect 494422 708982 530186 709218
rect 530422 708982 566186 709218
rect 566422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 8186 708598
rect 8422 708362 44186 708598
rect 44422 708362 80186 708598
rect 80422 708362 116186 708598
rect 116422 708362 152186 708598
rect 152422 708362 188186 708598
rect 188422 708362 224186 708598
rect 224422 708362 260186 708598
rect 260422 708362 296186 708598
rect 296422 708362 332186 708598
rect 332422 708362 368186 708598
rect 368422 708362 404186 708598
rect 404422 708362 440186 708598
rect 440422 708362 476186 708598
rect 476422 708362 512186 708598
rect 512422 708362 548186 708598
rect 548422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 8186 708278
rect 8422 708042 44186 708278
rect 44422 708042 80186 708278
rect 80422 708042 116186 708278
rect 116422 708042 152186 708278
rect 152422 708042 188186 708278
rect 188422 708042 224186 708278
rect 224422 708042 260186 708278
rect 260422 708042 296186 708278
rect 296422 708042 332186 708278
rect 332422 708042 368186 708278
rect 368422 708042 404186 708278
rect 404422 708042 440186 708278
rect 440422 708042 476186 708278
rect 476422 708042 512186 708278
rect 512422 708042 548186 708278
rect 548422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 22586 707658
rect 22822 707422 58586 707658
rect 58822 707422 94586 707658
rect 94822 707422 130586 707658
rect 130822 707422 166586 707658
rect 166822 707422 202586 707658
rect 202822 707422 238586 707658
rect 238822 707422 274586 707658
rect 274822 707422 310586 707658
rect 310822 707422 346586 707658
rect 346822 707422 382586 707658
rect 382822 707422 418586 707658
rect 418822 707422 454586 707658
rect 454822 707422 490586 707658
rect 490822 707422 526586 707658
rect 526822 707422 562586 707658
rect 562822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 22586 707338
rect 22822 707102 58586 707338
rect 58822 707102 94586 707338
rect 94822 707102 130586 707338
rect 130822 707102 166586 707338
rect 166822 707102 202586 707338
rect 202822 707102 238586 707338
rect 238822 707102 274586 707338
rect 274822 707102 310586 707338
rect 310822 707102 346586 707338
rect 346822 707102 382586 707338
rect 382822 707102 418586 707338
rect 418822 707102 454586 707338
rect 454822 707102 490586 707338
rect 490822 707102 526586 707338
rect 526822 707102 562586 707338
rect 562822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 4586 706718
rect 4822 706482 40586 706718
rect 40822 706482 76586 706718
rect 76822 706482 112586 706718
rect 112822 706482 148586 706718
rect 148822 706482 184586 706718
rect 184822 706482 220586 706718
rect 220822 706482 256586 706718
rect 256822 706482 292586 706718
rect 292822 706482 328586 706718
rect 328822 706482 364586 706718
rect 364822 706482 400586 706718
rect 400822 706482 436586 706718
rect 436822 706482 472586 706718
rect 472822 706482 508586 706718
rect 508822 706482 544586 706718
rect 544822 706482 580586 706718
rect 580822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 4586 706398
rect 4822 706162 40586 706398
rect 40822 706162 76586 706398
rect 76822 706162 112586 706398
rect 112822 706162 148586 706398
rect 148822 706162 184586 706398
rect 184822 706162 220586 706398
rect 220822 706162 256586 706398
rect 256822 706162 292586 706398
rect 292822 706162 328586 706398
rect 328822 706162 364586 706398
rect 364822 706162 400586 706398
rect 400822 706162 436586 706398
rect 436822 706162 472586 706398
rect 472822 706162 508586 706398
rect 508822 706162 544586 706398
rect 544822 706162 580586 706398
rect 580822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7636 697276 -7036 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590960 697276 591560 697278
rect -8576 697254 592500 697276
rect -8576 697018 -7454 697254
rect -7218 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591142 697254
rect 591378 697018 592500 697254
rect -8576 696934 592500 697018
rect -8576 696698 -7454 696934
rect -7218 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591142 696934
rect 591378 696698 592500 696934
rect -8576 696676 592500 696698
rect -7636 696674 -7036 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590960 696674 591560 696676
rect -5756 693676 -5156 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589080 693676 589680 693678
rect -6696 693654 590620 693676
rect -6696 693418 -5574 693654
rect -5338 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589262 693654
rect 589498 693418 590620 693654
rect -6696 693334 590620 693418
rect -6696 693098 -5574 693334
rect -5338 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589262 693334
rect 589498 693098 590620 693334
rect -6696 693076 590620 693098
rect -5756 693074 -5156 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589080 693074 589680 693076
rect -3876 690076 -3276 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587200 690076 587800 690078
rect -4816 690054 588740 690076
rect -4816 689818 -3694 690054
rect -3458 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587382 690054
rect 587618 689818 588740 690054
rect -4816 689734 588740 689818
rect -4816 689498 -3694 689734
rect -3458 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587382 689734
rect 587618 689498 588740 689734
rect -4816 689476 588740 689498
rect -3876 689474 -3276 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587200 689474 587800 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8576 679276 -7976 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591900 679276 592500 679278
rect -8576 679254 592500 679276
rect -8576 679018 -8394 679254
rect -8158 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 592082 679254
rect 592318 679018 592500 679254
rect -8576 678934 592500 679018
rect -8576 678698 -8394 678934
rect -8158 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 592082 678934
rect 592318 678698 592500 678934
rect -8576 678676 592500 678698
rect -8576 678674 -7976 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591900 678674 592500 678676
rect -6696 675676 -6096 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 590020 675676 590620 675678
rect -6696 675654 590620 675676
rect -6696 675418 -6514 675654
rect -6278 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590202 675654
rect 590438 675418 590620 675654
rect -6696 675334 590620 675418
rect -6696 675098 -6514 675334
rect -6278 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590202 675334
rect 590438 675098 590620 675334
rect -6696 675076 590620 675098
rect -6696 675074 -6096 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 590020 675074 590620 675076
rect -4816 672076 -4216 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588140 672076 588740 672078
rect -4816 672054 588740 672076
rect -4816 671818 -4634 672054
rect -4398 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588322 672054
rect 588558 671818 588740 672054
rect -4816 671734 588740 671818
rect -4816 671498 -4634 671734
rect -4398 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588322 671734
rect 588558 671498 588740 671734
rect -4816 671476 588740 671498
rect -4816 671474 -4216 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588140 671474 588740 671476
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -7636 661276 -7036 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590960 661276 591560 661278
rect -8576 661254 592500 661276
rect -8576 661018 -7454 661254
rect -7218 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591142 661254
rect 591378 661018 592500 661254
rect -8576 660934 592500 661018
rect -8576 660698 -7454 660934
rect -7218 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591142 660934
rect 591378 660698 592500 660934
rect -8576 660676 592500 660698
rect -7636 660674 -7036 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590960 660674 591560 660676
rect -5756 657676 -5156 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589080 657676 589680 657678
rect -6696 657654 590620 657676
rect -6696 657418 -5574 657654
rect -5338 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589262 657654
rect 589498 657418 590620 657654
rect -6696 657334 590620 657418
rect -6696 657098 -5574 657334
rect -5338 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589262 657334
rect 589498 657098 590620 657334
rect -6696 657076 590620 657098
rect -5756 657074 -5156 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589080 657074 589680 657076
rect -3876 654076 -3276 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587200 654076 587800 654078
rect -4816 654054 588740 654076
rect -4816 653818 -3694 654054
rect -3458 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587382 654054
rect 587618 653818 588740 654054
rect -4816 653734 588740 653818
rect -4816 653498 -3694 653734
rect -3458 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587382 653734
rect 587618 653498 588740 653734
rect -4816 653476 588740 653498
rect -3876 653474 -3276 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587200 653474 587800 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8576 643276 -7976 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591900 643276 592500 643278
rect -8576 643254 592500 643276
rect -8576 643018 -8394 643254
rect -8158 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 592082 643254
rect 592318 643018 592500 643254
rect -8576 642934 592500 643018
rect -8576 642698 -8394 642934
rect -8158 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 592082 642934
rect 592318 642698 592500 642934
rect -8576 642676 592500 642698
rect -8576 642674 -7976 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591900 642674 592500 642676
rect -6696 639676 -6096 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 590020 639676 590620 639678
rect -6696 639654 590620 639676
rect -6696 639418 -6514 639654
rect -6278 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590202 639654
rect 590438 639418 590620 639654
rect -6696 639334 590620 639418
rect -6696 639098 -6514 639334
rect -6278 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590202 639334
rect 590438 639098 590620 639334
rect -6696 639076 590620 639098
rect -6696 639074 -6096 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 590020 639074 590620 639076
rect -4816 636076 -4216 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588140 636076 588740 636078
rect -4816 636054 588740 636076
rect -4816 635818 -4634 636054
rect -4398 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588322 636054
rect 588558 635818 588740 636054
rect -4816 635734 588740 635818
rect -4816 635498 -4634 635734
rect -4398 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588322 635734
rect 588558 635498 588740 635734
rect -4816 635476 588740 635498
rect -4816 635474 -4216 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588140 635474 588740 635476
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -7636 625276 -7036 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590960 625276 591560 625278
rect -8576 625254 592500 625276
rect -8576 625018 -7454 625254
rect -7218 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591142 625254
rect 591378 625018 592500 625254
rect -8576 624934 592500 625018
rect -8576 624698 -7454 624934
rect -7218 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591142 624934
rect 591378 624698 592500 624934
rect -8576 624676 592500 624698
rect -7636 624674 -7036 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590960 624674 591560 624676
rect -5756 621676 -5156 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589080 621676 589680 621678
rect -6696 621654 590620 621676
rect -6696 621418 -5574 621654
rect -5338 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589262 621654
rect 589498 621418 590620 621654
rect -6696 621334 590620 621418
rect -6696 621098 -5574 621334
rect -5338 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589262 621334
rect 589498 621098 590620 621334
rect -6696 621076 590620 621098
rect -5756 621074 -5156 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589080 621074 589680 621076
rect -3876 618076 -3276 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587200 618076 587800 618078
rect -4816 618054 588740 618076
rect -4816 617818 -3694 618054
rect -3458 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587382 618054
rect 587618 617818 588740 618054
rect -4816 617734 588740 617818
rect -4816 617498 -3694 617734
rect -3458 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587382 617734
rect 587618 617498 588740 617734
rect -4816 617476 588740 617498
rect -3876 617474 -3276 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587200 617474 587800 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8576 607276 -7976 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591900 607276 592500 607278
rect -8576 607254 592500 607276
rect -8576 607018 -8394 607254
rect -8158 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 592082 607254
rect 592318 607018 592500 607254
rect -8576 606934 592500 607018
rect -8576 606698 -8394 606934
rect -8158 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 592082 606934
rect 592318 606698 592500 606934
rect -8576 606676 592500 606698
rect -8576 606674 -7976 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591900 606674 592500 606676
rect -6696 603676 -6096 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 590020 603676 590620 603678
rect -6696 603654 590620 603676
rect -6696 603418 -6514 603654
rect -6278 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590202 603654
rect 590438 603418 590620 603654
rect -6696 603334 590620 603418
rect -6696 603098 -6514 603334
rect -6278 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590202 603334
rect 590438 603098 590620 603334
rect -6696 603076 590620 603098
rect -6696 603074 -6096 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 590020 603074 590620 603076
rect -4816 600076 -4216 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588140 600076 588740 600078
rect -4816 600054 588740 600076
rect -4816 599818 -4634 600054
rect -4398 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588322 600054
rect 588558 599818 588740 600054
rect -4816 599734 588740 599818
rect -4816 599498 -4634 599734
rect -4398 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588322 599734
rect 588558 599498 588740 599734
rect -4816 599476 588740 599498
rect -4816 599474 -4216 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588140 599474 588740 599476
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -7636 589276 -7036 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590960 589276 591560 589278
rect -8576 589254 592500 589276
rect -8576 589018 -7454 589254
rect -7218 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591142 589254
rect 591378 589018 592500 589254
rect -8576 588934 592500 589018
rect -8576 588698 -7454 588934
rect -7218 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591142 588934
rect 591378 588698 592500 588934
rect -8576 588676 592500 588698
rect -7636 588674 -7036 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590960 588674 591560 588676
rect -5756 585676 -5156 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589080 585676 589680 585678
rect -6696 585654 590620 585676
rect -6696 585418 -5574 585654
rect -5338 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589262 585654
rect 589498 585418 590620 585654
rect -6696 585334 590620 585418
rect -6696 585098 -5574 585334
rect -5338 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589262 585334
rect 589498 585098 590620 585334
rect -6696 585076 590620 585098
rect -5756 585074 -5156 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589080 585074 589680 585076
rect -3876 582076 -3276 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587200 582076 587800 582078
rect -4816 582054 588740 582076
rect -4816 581818 -3694 582054
rect -3458 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587382 582054
rect 587618 581818 588740 582054
rect -4816 581734 588740 581818
rect -4816 581498 -3694 581734
rect -3458 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587382 581734
rect 587618 581498 588740 581734
rect -4816 581476 588740 581498
rect -3876 581474 -3276 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587200 581474 587800 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8576 571276 -7976 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 317604 571276 318204 571278
rect 353604 571276 354204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591900 571276 592500 571278
rect -8576 571254 592500 571276
rect -8576 571018 -8394 571254
rect -8158 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 317786 571254
rect 318022 571018 353786 571254
rect 354022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 592082 571254
rect 592318 571018 592500 571254
rect -8576 570934 592500 571018
rect -8576 570698 -8394 570934
rect -8158 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 317786 570934
rect 318022 570698 353786 570934
rect 354022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 592082 570934
rect 592318 570698 592500 570934
rect -8576 570676 592500 570698
rect -8576 570674 -7976 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 317604 570674 318204 570676
rect 353604 570674 354204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591900 570674 592500 570676
rect -6696 567676 -6096 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 314004 567676 314604 567678
rect 350004 567676 350604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 590020 567676 590620 567678
rect -6696 567654 590620 567676
rect -6696 567418 -6514 567654
rect -6278 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 314186 567654
rect 314422 567418 350186 567654
rect 350422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590202 567654
rect 590438 567418 590620 567654
rect -6696 567334 590620 567418
rect -6696 567098 -6514 567334
rect -6278 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 314186 567334
rect 314422 567098 350186 567334
rect 350422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590202 567334
rect 590438 567098 590620 567334
rect -6696 567076 590620 567098
rect -6696 567074 -6096 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 314004 567074 314604 567076
rect 350004 567074 350604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 590020 567074 590620 567076
rect -4816 564076 -4216 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588140 564076 588740 564078
rect -4816 564054 588740 564076
rect -4816 563818 -4634 564054
rect -4398 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588322 564054
rect 588558 563818 588740 564054
rect -4816 563734 588740 563818
rect -4816 563498 -4634 563734
rect -4398 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588322 563734
rect 588558 563498 588740 563734
rect -4816 563476 588740 563498
rect -4816 563474 -4216 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588140 563474 588740 563476
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -7636 553276 -7036 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590960 553276 591560 553278
rect -8576 553254 592500 553276
rect -8576 553018 -7454 553254
rect -7218 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591142 553254
rect 591378 553018 592500 553254
rect -8576 552934 592500 553018
rect -8576 552698 -7454 552934
rect -7218 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591142 552934
rect 591378 552698 592500 552934
rect -8576 552676 592500 552698
rect -7636 552674 -7036 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590960 552674 591560 552676
rect -5756 549676 -5156 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589080 549676 589680 549678
rect -6696 549654 590620 549676
rect -6696 549418 -5574 549654
rect -5338 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589262 549654
rect 589498 549418 590620 549654
rect -6696 549334 590620 549418
rect -6696 549098 -5574 549334
rect -5338 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589262 549334
rect 589498 549098 590620 549334
rect -6696 549076 590620 549098
rect -5756 549074 -5156 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589080 549074 589680 549076
rect -3876 546076 -3276 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587200 546076 587800 546078
rect -4816 546054 588740 546076
rect -4816 545818 -3694 546054
rect -3458 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587382 546054
rect 587618 545818 588740 546054
rect -4816 545734 588740 545818
rect -4816 545498 -3694 545734
rect -3458 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587382 545734
rect 587618 545498 588740 545734
rect -4816 545476 588740 545498
rect -3876 545474 -3276 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587200 545474 587800 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8576 535276 -7976 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 101604 535276 102204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 209604 535276 210204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591900 535276 592500 535278
rect -8576 535254 592500 535276
rect -8576 535018 -8394 535254
rect -8158 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 101786 535254
rect 102022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 209786 535254
rect 210022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 592082 535254
rect 592318 535018 592500 535254
rect -8576 534934 592500 535018
rect -8576 534698 -8394 534934
rect -8158 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 101786 534934
rect 102022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 209786 534934
rect 210022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 592082 534934
rect 592318 534698 592500 534934
rect -8576 534676 592500 534698
rect -8576 534674 -7976 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 101604 534674 102204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 209604 534674 210204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591900 534674 592500 534676
rect -6696 531676 -6096 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 98004 531676 98604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 206004 531676 206604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 590020 531676 590620 531678
rect -6696 531654 590620 531676
rect -6696 531418 -6514 531654
rect -6278 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 98186 531654
rect 98422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 206186 531654
rect 206422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590202 531654
rect 590438 531418 590620 531654
rect -6696 531334 590620 531418
rect -6696 531098 -6514 531334
rect -6278 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 98186 531334
rect 98422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 206186 531334
rect 206422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590202 531334
rect 590438 531098 590620 531334
rect -6696 531076 590620 531098
rect -6696 531074 -6096 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 98004 531074 98604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 206004 531074 206604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 590020 531074 590620 531076
rect -4816 528076 -4216 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588140 528076 588740 528078
rect -4816 528054 588740 528076
rect -4816 527818 -4634 528054
rect -4398 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588322 528054
rect 588558 527818 588740 528054
rect -4816 527734 588740 527818
rect -4816 527498 -4634 527734
rect -4398 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588322 527734
rect 588558 527498 588740 527734
rect -4816 527476 588740 527498
rect -4816 527474 -4216 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588140 527474 588740 527476
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586260 523874 586860 523876
rect -7636 517276 -7036 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 299604 517276 300204 517278
rect 335604 517276 336204 517278
rect 371604 517276 372204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590960 517276 591560 517278
rect -8576 517254 592500 517276
rect -8576 517018 -7454 517254
rect -7218 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 299786 517254
rect 300022 517018 335786 517254
rect 336022 517018 371786 517254
rect 372022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591142 517254
rect 591378 517018 592500 517254
rect -8576 516934 592500 517018
rect -8576 516698 -7454 516934
rect -7218 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 299786 516934
rect 300022 516698 335786 516934
rect 336022 516698 371786 516934
rect 372022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591142 516934
rect 591378 516698 592500 516934
rect -8576 516676 592500 516698
rect -7636 516674 -7036 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 299604 516674 300204 516676
rect 335604 516674 336204 516676
rect 371604 516674 372204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590960 516674 591560 516676
rect -5756 513676 -5156 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589080 513676 589680 513678
rect -6696 513654 590620 513676
rect -6696 513418 -5574 513654
rect -5338 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589262 513654
rect 589498 513418 590620 513654
rect -6696 513334 590620 513418
rect -6696 513098 -5574 513334
rect -5338 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589262 513334
rect 589498 513098 590620 513334
rect -6696 513076 590620 513098
rect -5756 513074 -5156 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589080 513074 589680 513076
rect -3876 510076 -3276 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587200 510076 587800 510078
rect -4816 510054 588740 510076
rect -4816 509818 -3694 510054
rect -3458 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587382 510054
rect 587618 509818 588740 510054
rect -4816 509734 588740 509818
rect -4816 509498 -3694 509734
rect -3458 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587382 509734
rect 587618 509498 588740 509734
rect -4816 509476 588740 509498
rect -3876 509474 -3276 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587200 509474 587800 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8576 499276 -7976 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591900 499276 592500 499278
rect -8576 499254 592500 499276
rect -8576 499018 -8394 499254
rect -8158 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 592082 499254
rect 592318 499018 592500 499254
rect -8576 498934 592500 499018
rect -8576 498698 -8394 498934
rect -8158 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 592082 498934
rect 592318 498698 592500 498934
rect -8576 498676 592500 498698
rect -8576 498674 -7976 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591900 498674 592500 498676
rect -6696 495676 -6096 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 590020 495676 590620 495678
rect -6696 495654 590620 495676
rect -6696 495418 -6514 495654
rect -6278 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590202 495654
rect 590438 495418 590620 495654
rect -6696 495334 590620 495418
rect -6696 495098 -6514 495334
rect -6278 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590202 495334
rect 590438 495098 590620 495334
rect -6696 495076 590620 495098
rect -6696 495074 -6096 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 590020 495074 590620 495076
rect -4816 492076 -4216 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588140 492076 588740 492078
rect -4816 492054 588740 492076
rect -4816 491818 -4634 492054
rect -4398 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588322 492054
rect 588558 491818 588740 492054
rect -4816 491734 588740 491818
rect -4816 491498 -4634 491734
rect -4398 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588322 491734
rect 588558 491498 588740 491734
rect -4816 491476 588740 491498
rect -4816 491474 -4216 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588140 491474 588740 491476
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -7636 481276 -7036 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 263604 481276 264204 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590960 481276 591560 481278
rect -8576 481254 592500 481276
rect -8576 481018 -7454 481254
rect -7218 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 263786 481254
rect 264022 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591142 481254
rect 591378 481018 592500 481254
rect -8576 480934 592500 481018
rect -8576 480698 -7454 480934
rect -7218 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 263786 480934
rect 264022 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591142 480934
rect 591378 480698 592500 480934
rect -8576 480676 592500 480698
rect -7636 480674 -7036 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 263604 480674 264204 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590960 480674 591560 480676
rect -5756 477676 -5156 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 260004 477676 260604 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589080 477676 589680 477678
rect -6696 477654 590620 477676
rect -6696 477418 -5574 477654
rect -5338 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 260186 477654
rect 260422 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589262 477654
rect 589498 477418 590620 477654
rect -6696 477334 590620 477418
rect -6696 477098 -5574 477334
rect -5338 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 260186 477334
rect 260422 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589262 477334
rect 589498 477098 590620 477334
rect -6696 477076 590620 477098
rect -5756 477074 -5156 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 260004 477074 260604 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589080 477074 589680 477076
rect -3876 474076 -3276 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587200 474076 587800 474078
rect -4816 474054 588740 474076
rect -4816 473818 -3694 474054
rect -3458 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587382 474054
rect 587618 473818 588740 474054
rect -4816 473734 588740 473818
rect -4816 473498 -3694 473734
rect -3458 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587382 473734
rect 587618 473498 588740 473734
rect -4816 473476 588740 473498
rect -3876 473474 -3276 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587200 473474 587800 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8576 463276 -7976 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 281604 463276 282204 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591900 463276 592500 463278
rect -8576 463254 592500 463276
rect -8576 463018 -8394 463254
rect -8158 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 281786 463254
rect 282022 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 592082 463254
rect 592318 463018 592500 463254
rect -8576 462934 592500 463018
rect -8576 462698 -8394 462934
rect -8158 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 281786 462934
rect 282022 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 592082 462934
rect 592318 462698 592500 462934
rect -8576 462676 592500 462698
rect -8576 462674 -7976 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 281604 462674 282204 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591900 462674 592500 462676
rect -6696 459676 -6096 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 278004 459676 278604 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 590020 459676 590620 459678
rect -6696 459654 590620 459676
rect -6696 459418 -6514 459654
rect -6278 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 278186 459654
rect 278422 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590202 459654
rect 590438 459418 590620 459654
rect -6696 459334 590620 459418
rect -6696 459098 -6514 459334
rect -6278 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 278186 459334
rect 278422 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590202 459334
rect 590438 459098 590620 459334
rect -6696 459076 590620 459098
rect -6696 459074 -6096 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 278004 459074 278604 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 590020 459074 590620 459076
rect -4816 456076 -4216 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588140 456076 588740 456078
rect -4816 456054 588740 456076
rect -4816 455818 -4634 456054
rect -4398 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588322 456054
rect 588558 455818 588740 456054
rect -4816 455734 588740 455818
rect -4816 455498 -4634 455734
rect -4398 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588322 455734
rect 588558 455498 588740 455734
rect -4816 455476 588740 455498
rect -4816 455474 -4216 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588140 455474 588740 455476
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -7636 445276 -7036 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590960 445276 591560 445278
rect -8576 445254 592500 445276
rect -8576 445018 -7454 445254
rect -7218 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591142 445254
rect 591378 445018 592500 445254
rect -8576 444934 592500 445018
rect -8576 444698 -7454 444934
rect -7218 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591142 444934
rect 591378 444698 592500 444934
rect -8576 444676 592500 444698
rect -7636 444674 -7036 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590960 444674 591560 444676
rect -5756 441676 -5156 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 260004 441676 260604 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589080 441676 589680 441678
rect -6696 441654 590620 441676
rect -6696 441418 -5574 441654
rect -5338 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 260186 441654
rect 260422 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589262 441654
rect 589498 441418 590620 441654
rect -6696 441334 590620 441418
rect -6696 441098 -5574 441334
rect -5338 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 260186 441334
rect 260422 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589262 441334
rect 589498 441098 590620 441334
rect -6696 441076 590620 441098
rect -5756 441074 -5156 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 260004 441074 260604 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589080 441074 589680 441076
rect -3876 438076 -3276 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587200 438076 587800 438078
rect -4816 438054 588740 438076
rect -4816 437818 -3694 438054
rect -3458 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587382 438054
rect 587618 437818 588740 438054
rect -4816 437734 588740 437818
rect -4816 437498 -3694 437734
rect -3458 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587382 437734
rect 587618 437498 588740 437734
rect -4816 437476 588740 437498
rect -3876 437474 -3276 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587200 437474 587800 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8576 427276 -7976 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 281604 427276 282204 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591900 427276 592500 427278
rect -8576 427254 592500 427276
rect -8576 427018 -8394 427254
rect -8158 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 281786 427254
rect 282022 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 592082 427254
rect 592318 427018 592500 427254
rect -8576 426934 592500 427018
rect -8576 426698 -8394 426934
rect -8158 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 281786 426934
rect 282022 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 592082 426934
rect 592318 426698 592500 426934
rect -8576 426676 592500 426698
rect -8576 426674 -7976 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 281604 426674 282204 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591900 426674 592500 426676
rect -6696 423676 -6096 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 278004 423676 278604 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 590020 423676 590620 423678
rect -6696 423654 590620 423676
rect -6696 423418 -6514 423654
rect -6278 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 278186 423654
rect 278422 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590202 423654
rect 590438 423418 590620 423654
rect -6696 423334 590620 423418
rect -6696 423098 -6514 423334
rect -6278 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 278186 423334
rect 278422 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590202 423334
rect 590438 423098 590620 423334
rect -6696 423076 590620 423098
rect -6696 423074 -6096 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 278004 423074 278604 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 590020 423074 590620 423076
rect -4816 420076 -4216 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 238404 420076 239004 420078
rect 274404 420076 275004 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588140 420076 588740 420078
rect -4816 420054 588740 420076
rect -4816 419818 -4634 420054
rect -4398 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 238586 420054
rect 238822 419818 274586 420054
rect 274822 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588322 420054
rect 588558 419818 588740 420054
rect -4816 419734 588740 419818
rect -4816 419498 -4634 419734
rect -4398 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 238586 419734
rect 238822 419498 274586 419734
rect 274822 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588322 419734
rect 588558 419498 588740 419734
rect -4816 419476 588740 419498
rect -4816 419474 -4216 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 238404 419474 239004 419476
rect 274404 419474 275004 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588140 419474 588740 419476
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect -7636 409276 -7036 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590960 409276 591560 409278
rect -8576 409254 592500 409276
rect -8576 409018 -7454 409254
rect -7218 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591142 409254
rect 591378 409018 592500 409254
rect -8576 408934 592500 409018
rect -8576 408698 -7454 408934
rect -7218 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591142 408934
rect 591378 408698 592500 408934
rect -8576 408676 592500 408698
rect -7636 408674 -7036 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590960 408674 591560 408676
rect -5756 405676 -5156 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589080 405676 589680 405678
rect -6696 405654 590620 405676
rect -6696 405418 -5574 405654
rect -5338 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589262 405654
rect 589498 405418 590620 405654
rect -6696 405334 590620 405418
rect -6696 405098 -5574 405334
rect -5338 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589262 405334
rect 589498 405098 590620 405334
rect -6696 405076 590620 405098
rect -5756 405074 -5156 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589080 405074 589680 405076
rect -3876 402076 -3276 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587200 402076 587800 402078
rect -4816 402054 588740 402076
rect -4816 401818 -3694 402054
rect -3458 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587382 402054
rect 587618 401818 588740 402054
rect -4816 401734 588740 401818
rect -4816 401498 -3694 401734
rect -3458 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587382 401734
rect 587618 401498 588740 401734
rect -4816 401476 588740 401498
rect -3876 401474 -3276 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587200 401474 587800 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8576 391276 -7976 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 101604 391276 102204 391278
rect 137604 391276 138204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591900 391276 592500 391278
rect -8576 391254 592500 391276
rect -8576 391018 -8394 391254
rect -8158 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 101786 391254
rect 102022 391018 137786 391254
rect 138022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 592082 391254
rect 592318 391018 592500 391254
rect -8576 390934 592500 391018
rect -8576 390698 -8394 390934
rect -8158 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 101786 390934
rect 102022 390698 137786 390934
rect 138022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 592082 390934
rect 592318 390698 592500 390934
rect -8576 390676 592500 390698
rect -8576 390674 -7976 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 101604 390674 102204 390676
rect 137604 390674 138204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591900 390674 592500 390676
rect -6696 387676 -6096 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 98004 387676 98604 387678
rect 134004 387676 134604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 590020 387676 590620 387678
rect -6696 387654 590620 387676
rect -6696 387418 -6514 387654
rect -6278 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 98186 387654
rect 98422 387418 134186 387654
rect 134422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590202 387654
rect 590438 387418 590620 387654
rect -6696 387334 590620 387418
rect -6696 387098 -6514 387334
rect -6278 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 98186 387334
rect 98422 387098 134186 387334
rect 134422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590202 387334
rect 590438 387098 590620 387334
rect -6696 387076 590620 387098
rect -6696 387074 -6096 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 98004 387074 98604 387076
rect 134004 387074 134604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 590020 387074 590620 387076
rect -4816 384076 -4216 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588140 384076 588740 384078
rect -4816 384054 588740 384076
rect -4816 383818 -4634 384054
rect -4398 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588322 384054
rect 588558 383818 588740 384054
rect -4816 383734 588740 383818
rect -4816 383498 -4634 383734
rect -4398 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588322 383734
rect 588558 383498 588740 383734
rect -4816 383476 588740 383498
rect -4816 383474 -4216 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588140 383474 588740 383476
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -7636 373276 -7036 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 83604 373276 84204 373278
rect 119604 373276 120204 373278
rect 407604 373276 408204 373278
rect 443604 373276 444204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590960 373276 591560 373278
rect -8576 373254 592500 373276
rect -8576 373018 -7454 373254
rect -7218 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 83786 373254
rect 84022 373018 119786 373254
rect 120022 373018 407786 373254
rect 408022 373018 443786 373254
rect 444022 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591142 373254
rect 591378 373018 592500 373254
rect -8576 372934 592500 373018
rect -8576 372698 -7454 372934
rect -7218 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 83786 372934
rect 84022 372698 119786 372934
rect 120022 372698 407786 372934
rect 408022 372698 443786 372934
rect 444022 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591142 372934
rect 591378 372698 592500 372934
rect -8576 372676 592500 372698
rect -7636 372674 -7036 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 83604 372674 84204 372676
rect 119604 372674 120204 372676
rect 407604 372674 408204 372676
rect 443604 372674 444204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590960 372674 591560 372676
rect -5756 369676 -5156 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 116004 369676 116604 369678
rect 152004 369676 152604 369678
rect 404004 369676 404604 369678
rect 440004 369676 440604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589080 369676 589680 369678
rect -6696 369654 590620 369676
rect -6696 369418 -5574 369654
rect -5338 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 116186 369654
rect 116422 369418 152186 369654
rect 152422 369418 404186 369654
rect 404422 369418 440186 369654
rect 440422 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589262 369654
rect 589498 369418 590620 369654
rect -6696 369334 590620 369418
rect -6696 369098 -5574 369334
rect -5338 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 116186 369334
rect 116422 369098 152186 369334
rect 152422 369098 404186 369334
rect 404422 369098 440186 369334
rect 440422 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589262 369334
rect 589498 369098 590620 369334
rect -6696 369076 590620 369098
rect -5756 369074 -5156 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 116004 369074 116604 369076
rect 152004 369074 152604 369076
rect 404004 369074 404604 369076
rect 440004 369074 440604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589080 369074 589680 369076
rect -3876 366076 -3276 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 148404 366076 149004 366078
rect 400404 366076 401004 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587200 366076 587800 366078
rect -4816 366054 588740 366076
rect -4816 365818 -3694 366054
rect -3458 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 148586 366054
rect 148822 365818 400586 366054
rect 400822 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587382 366054
rect 587618 365818 588740 366054
rect -4816 365734 588740 365818
rect -4816 365498 -3694 365734
rect -3458 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 148586 365734
rect 148822 365498 400586 365734
rect 400822 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587382 365734
rect 587618 365498 588740 365734
rect -4816 365476 588740 365498
rect -3876 365474 -3276 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 148404 365474 149004 365476
rect 400404 365474 401004 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587200 365474 587800 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8576 355276 -7976 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 101604 355276 102204 355278
rect 137604 355276 138204 355278
rect 425604 355276 426204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591900 355276 592500 355278
rect -8576 355254 592500 355276
rect -8576 355018 -8394 355254
rect -8158 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 101786 355254
rect 102022 355018 137786 355254
rect 138022 355018 425786 355254
rect 426022 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 592082 355254
rect 592318 355018 592500 355254
rect -8576 354934 592500 355018
rect -8576 354698 -8394 354934
rect -8158 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 101786 354934
rect 102022 354698 137786 354934
rect 138022 354698 425786 354934
rect 426022 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 592082 354934
rect 592318 354698 592500 354934
rect -8576 354676 592500 354698
rect -8576 354674 -7976 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 101604 354674 102204 354676
rect 137604 354674 138204 354676
rect 425604 354674 426204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591900 354674 592500 354676
rect -6696 351676 -6096 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 98004 351676 98604 351678
rect 134004 351676 134604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 590020 351676 590620 351678
rect -6696 351654 590620 351676
rect -6696 351418 -6514 351654
rect -6278 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 98186 351654
rect 98422 351418 134186 351654
rect 134422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590202 351654
rect 590438 351418 590620 351654
rect -6696 351334 590620 351418
rect -6696 351098 -6514 351334
rect -6278 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 98186 351334
rect 98422 351098 134186 351334
rect 134422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590202 351334
rect 590438 351098 590620 351334
rect -6696 351076 590620 351098
rect -6696 351074 -6096 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 98004 351074 98604 351076
rect 134004 351074 134604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 590020 351074 590620 351076
rect -4816 348076 -4216 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588140 348076 588740 348078
rect -4816 348054 588740 348076
rect -4816 347818 -4634 348054
rect -4398 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588322 348054
rect 588558 347818 588740 348054
rect -4816 347734 588740 347818
rect -4816 347498 -4634 347734
rect -4398 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588322 347734
rect 588558 347498 588740 347734
rect -4816 347476 588740 347498
rect -4816 347474 -4216 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588140 347474 588740 347476
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -7636 337276 -7036 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 407604 337276 408204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590960 337276 591560 337278
rect -8576 337254 592500 337276
rect -8576 337018 -7454 337254
rect -7218 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 407786 337254
rect 408022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591142 337254
rect 591378 337018 592500 337254
rect -8576 336934 592500 337018
rect -8576 336698 -7454 336934
rect -7218 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 407786 336934
rect 408022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591142 336934
rect 591378 336698 592500 336934
rect -8576 336676 592500 336698
rect -7636 336674 -7036 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 407604 336674 408204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590960 336674 591560 336676
rect -5756 333676 -5156 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 404004 333676 404604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589080 333676 589680 333678
rect -6696 333654 590620 333676
rect -6696 333418 -5574 333654
rect -5338 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 404186 333654
rect 404422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589262 333654
rect 589498 333418 590620 333654
rect -6696 333334 590620 333418
rect -6696 333098 -5574 333334
rect -5338 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 404186 333334
rect 404422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589262 333334
rect 589498 333098 590620 333334
rect -6696 333076 590620 333098
rect -5756 333074 -5156 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 404004 333074 404604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589080 333074 589680 333076
rect -3876 330076 -3276 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587200 330076 587800 330078
rect -4816 330054 588740 330076
rect -4816 329818 -3694 330054
rect -3458 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587382 330054
rect 587618 329818 588740 330054
rect -4816 329734 588740 329818
rect -4816 329498 -3694 329734
rect -3458 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587382 329734
rect 587618 329498 588740 329734
rect -4816 329476 588740 329498
rect -3876 329474 -3276 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587200 329474 587800 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8576 319276 -7976 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591900 319276 592500 319278
rect -8576 319254 592500 319276
rect -8576 319018 -8394 319254
rect -8158 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 592082 319254
rect 592318 319018 592500 319254
rect -8576 318934 592500 319018
rect -8576 318698 -8394 318934
rect -8158 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 592082 318934
rect 592318 318698 592500 318934
rect -8576 318676 592500 318698
rect -8576 318674 -7976 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591900 318674 592500 318676
rect -6696 315676 -6096 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 590020 315676 590620 315678
rect -6696 315654 590620 315676
rect -6696 315418 -6514 315654
rect -6278 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590202 315654
rect 590438 315418 590620 315654
rect -6696 315334 590620 315418
rect -6696 315098 -6514 315334
rect -6278 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590202 315334
rect 590438 315098 590620 315334
rect -6696 315076 590620 315098
rect -6696 315074 -6096 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 590020 315074 590620 315076
rect -4816 312076 -4216 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588140 312076 588740 312078
rect -4816 312054 588740 312076
rect -4816 311818 -4634 312054
rect -4398 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588322 312054
rect 588558 311818 588740 312054
rect -4816 311734 588740 311818
rect -4816 311498 -4634 311734
rect -4398 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588322 311734
rect 588558 311498 588740 311734
rect -4816 311476 588740 311498
rect -4816 311474 -4216 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588140 311474 588740 311476
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -7636 301276 -7036 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590960 301276 591560 301278
rect -8576 301254 592500 301276
rect -8576 301018 -7454 301254
rect -7218 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591142 301254
rect 591378 301018 592500 301254
rect -8576 300934 592500 301018
rect -8576 300698 -7454 300934
rect -7218 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591142 300934
rect 591378 300698 592500 300934
rect -8576 300676 592500 300698
rect -7636 300674 -7036 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590960 300674 591560 300676
rect -5756 297676 -5156 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589080 297676 589680 297678
rect -6696 297654 590620 297676
rect -6696 297418 -5574 297654
rect -5338 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589262 297654
rect 589498 297418 590620 297654
rect -6696 297334 590620 297418
rect -6696 297098 -5574 297334
rect -5338 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589262 297334
rect 589498 297098 590620 297334
rect -6696 297076 590620 297098
rect -5756 297074 -5156 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589080 297074 589680 297076
rect -3876 294076 -3276 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587200 294076 587800 294078
rect -4816 294054 588740 294076
rect -4816 293818 -3694 294054
rect -3458 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587382 294054
rect 587618 293818 588740 294054
rect -4816 293734 588740 293818
rect -4816 293498 -3694 293734
rect -3458 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587382 293734
rect 587618 293498 588740 293734
rect -4816 293476 588740 293498
rect -3876 293474 -3276 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587200 293474 587800 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8576 283276 -7976 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591900 283276 592500 283278
rect -8576 283254 592500 283276
rect -8576 283018 -8394 283254
rect -8158 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 592082 283254
rect 592318 283018 592500 283254
rect -8576 282934 592500 283018
rect -8576 282698 -8394 282934
rect -8158 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 592082 282934
rect 592318 282698 592500 282934
rect -8576 282676 592500 282698
rect -8576 282674 -7976 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591900 282674 592500 282676
rect -6696 279676 -6096 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 590020 279676 590620 279678
rect -6696 279654 590620 279676
rect -6696 279418 -6514 279654
rect -6278 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590202 279654
rect 590438 279418 590620 279654
rect -6696 279334 590620 279418
rect -6696 279098 -6514 279334
rect -6278 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590202 279334
rect 590438 279098 590620 279334
rect -6696 279076 590620 279098
rect -6696 279074 -6096 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 590020 279074 590620 279076
rect -4816 276076 -4216 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588140 276076 588740 276078
rect -4816 276054 588740 276076
rect -4816 275818 -4634 276054
rect -4398 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588322 276054
rect 588558 275818 588740 276054
rect -4816 275734 588740 275818
rect -4816 275498 -4634 275734
rect -4398 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588322 275734
rect 588558 275498 588740 275734
rect -4816 275476 588740 275498
rect -4816 275474 -4216 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588140 275474 588740 275476
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -7636 265276 -7036 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590960 265276 591560 265278
rect -8576 265254 592500 265276
rect -8576 265018 -7454 265254
rect -7218 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591142 265254
rect 591378 265018 592500 265254
rect -8576 264934 592500 265018
rect -8576 264698 -7454 264934
rect -7218 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591142 264934
rect 591378 264698 592500 264934
rect -8576 264676 592500 264698
rect -7636 264674 -7036 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590960 264674 591560 264676
rect -5756 261676 -5156 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589080 261676 589680 261678
rect -6696 261654 590620 261676
rect -6696 261418 -5574 261654
rect -5338 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589262 261654
rect 589498 261418 590620 261654
rect -6696 261334 590620 261418
rect -6696 261098 -5574 261334
rect -5338 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589262 261334
rect 589498 261098 590620 261334
rect -6696 261076 590620 261098
rect -5756 261074 -5156 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589080 261074 589680 261076
rect -3876 258076 -3276 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587200 258076 587800 258078
rect -4816 258054 588740 258076
rect -4816 257818 -3694 258054
rect -3458 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587382 258054
rect 587618 257818 588740 258054
rect -4816 257734 588740 257818
rect -4816 257498 -3694 257734
rect -3458 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587382 257734
rect 587618 257498 588740 257734
rect -4816 257476 588740 257498
rect -3876 257474 -3276 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587200 257474 587800 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8576 247276 -7976 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591900 247276 592500 247278
rect -8576 247254 592500 247276
rect -8576 247018 -8394 247254
rect -8158 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 592082 247254
rect 592318 247018 592500 247254
rect -8576 246934 592500 247018
rect -8576 246698 -8394 246934
rect -8158 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 592082 246934
rect 592318 246698 592500 246934
rect -8576 246676 592500 246698
rect -8576 246674 -7976 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591900 246674 592500 246676
rect -6696 243676 -6096 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 590020 243676 590620 243678
rect -6696 243654 590620 243676
rect -6696 243418 -6514 243654
rect -6278 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590202 243654
rect 590438 243418 590620 243654
rect -6696 243334 590620 243418
rect -6696 243098 -6514 243334
rect -6278 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590202 243334
rect 590438 243098 590620 243334
rect -6696 243076 590620 243098
rect -6696 243074 -6096 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 590020 243074 590620 243076
rect -4816 240076 -4216 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588140 240076 588740 240078
rect -4816 240054 588740 240076
rect -4816 239818 -4634 240054
rect -4398 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588322 240054
rect 588558 239818 588740 240054
rect -4816 239734 588740 239818
rect -4816 239498 -4634 239734
rect -4398 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588322 239734
rect 588558 239498 588740 239734
rect -4816 239476 588740 239498
rect -4816 239474 -4216 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588140 239474 588740 239476
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -7636 229276 -7036 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590960 229276 591560 229278
rect -8576 229254 592500 229276
rect -8576 229018 -7454 229254
rect -7218 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591142 229254
rect 591378 229018 592500 229254
rect -8576 228934 592500 229018
rect -8576 228698 -7454 228934
rect -7218 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591142 228934
rect 591378 228698 592500 228934
rect -8576 228676 592500 228698
rect -7636 228674 -7036 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590960 228674 591560 228676
rect -5756 225676 -5156 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589080 225676 589680 225678
rect -6696 225654 590620 225676
rect -6696 225418 -5574 225654
rect -5338 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589262 225654
rect 589498 225418 590620 225654
rect -6696 225334 590620 225418
rect -6696 225098 -5574 225334
rect -5338 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589262 225334
rect 589498 225098 590620 225334
rect -6696 225076 590620 225098
rect -5756 225074 -5156 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589080 225074 589680 225076
rect -3876 222076 -3276 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587200 222076 587800 222078
rect -4816 222054 588740 222076
rect -4816 221818 -3694 222054
rect -3458 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587382 222054
rect 587618 221818 588740 222054
rect -4816 221734 588740 221818
rect -4816 221498 -3694 221734
rect -3458 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587382 221734
rect 587618 221498 588740 221734
rect -4816 221476 588740 221498
rect -3876 221474 -3276 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587200 221474 587800 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8576 211276 -7976 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591900 211276 592500 211278
rect -8576 211254 592500 211276
rect -8576 211018 -8394 211254
rect -8158 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 592082 211254
rect 592318 211018 592500 211254
rect -8576 210934 592500 211018
rect -8576 210698 -8394 210934
rect -8158 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 592082 210934
rect 592318 210698 592500 210934
rect -8576 210676 592500 210698
rect -8576 210674 -7976 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591900 210674 592500 210676
rect -6696 207676 -6096 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 590020 207676 590620 207678
rect -6696 207654 590620 207676
rect -6696 207418 -6514 207654
rect -6278 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590202 207654
rect 590438 207418 590620 207654
rect -6696 207334 590620 207418
rect -6696 207098 -6514 207334
rect -6278 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590202 207334
rect 590438 207098 590620 207334
rect -6696 207076 590620 207098
rect -6696 207074 -6096 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 590020 207074 590620 207076
rect -4816 204076 -4216 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588140 204076 588740 204078
rect -4816 204054 588740 204076
rect -4816 203818 -4634 204054
rect -4398 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588322 204054
rect 588558 203818 588740 204054
rect -4816 203734 588740 203818
rect -4816 203498 -4634 203734
rect -4398 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588322 203734
rect 588558 203498 588740 203734
rect -4816 203476 588740 203498
rect -4816 203474 -4216 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588140 203474 588740 203476
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -7636 193276 -7036 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590960 193276 591560 193278
rect -8576 193254 592500 193276
rect -8576 193018 -7454 193254
rect -7218 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591142 193254
rect 591378 193018 592500 193254
rect -8576 192934 592500 193018
rect -8576 192698 -7454 192934
rect -7218 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591142 192934
rect 591378 192698 592500 192934
rect -8576 192676 592500 192698
rect -7636 192674 -7036 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590960 192674 591560 192676
rect -5756 189676 -5156 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589080 189676 589680 189678
rect -6696 189654 590620 189676
rect -6696 189418 -5574 189654
rect -5338 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589262 189654
rect 589498 189418 590620 189654
rect -6696 189334 590620 189418
rect -6696 189098 -5574 189334
rect -5338 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589262 189334
rect 589498 189098 590620 189334
rect -6696 189076 590620 189098
rect -5756 189074 -5156 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589080 189074 589680 189076
rect -3876 186076 -3276 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587200 186076 587800 186078
rect -4816 186054 588740 186076
rect -4816 185818 -3694 186054
rect -3458 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587382 186054
rect 587618 185818 588740 186054
rect -4816 185734 588740 185818
rect -4816 185498 -3694 185734
rect -3458 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587382 185734
rect 587618 185498 588740 185734
rect -4816 185476 588740 185498
rect -3876 185474 -3276 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587200 185474 587800 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8576 175276 -7976 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591900 175276 592500 175278
rect -8576 175254 592500 175276
rect -8576 175018 -8394 175254
rect -8158 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 592082 175254
rect 592318 175018 592500 175254
rect -8576 174934 592500 175018
rect -8576 174698 -8394 174934
rect -8158 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 592082 174934
rect 592318 174698 592500 174934
rect -8576 174676 592500 174698
rect -8576 174674 -7976 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591900 174674 592500 174676
rect -6696 171676 -6096 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 590020 171676 590620 171678
rect -6696 171654 590620 171676
rect -6696 171418 -6514 171654
rect -6278 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590202 171654
rect 590438 171418 590620 171654
rect -6696 171334 590620 171418
rect -6696 171098 -6514 171334
rect -6278 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590202 171334
rect 590438 171098 590620 171334
rect -6696 171076 590620 171098
rect -6696 171074 -6096 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 590020 171074 590620 171076
rect -4816 168076 -4216 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588140 168076 588740 168078
rect -4816 168054 588740 168076
rect -4816 167818 -4634 168054
rect -4398 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588322 168054
rect 588558 167818 588740 168054
rect -4816 167734 588740 167818
rect -4816 167498 -4634 167734
rect -4398 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588322 167734
rect 588558 167498 588740 167734
rect -4816 167476 588740 167498
rect -4816 167474 -4216 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588140 167474 588740 167476
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -7636 157276 -7036 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590960 157276 591560 157278
rect -8576 157254 592500 157276
rect -8576 157018 -7454 157254
rect -7218 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591142 157254
rect 591378 157018 592500 157254
rect -8576 156934 592500 157018
rect -8576 156698 -7454 156934
rect -7218 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591142 156934
rect 591378 156698 592500 156934
rect -8576 156676 592500 156698
rect -7636 156674 -7036 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590960 156674 591560 156676
rect -5756 153676 -5156 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589080 153676 589680 153678
rect -6696 153654 590620 153676
rect -6696 153418 -5574 153654
rect -5338 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589262 153654
rect 589498 153418 590620 153654
rect -6696 153334 590620 153418
rect -6696 153098 -5574 153334
rect -5338 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589262 153334
rect 589498 153098 590620 153334
rect -6696 153076 590620 153098
rect -5756 153074 -5156 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589080 153074 589680 153076
rect -3876 150076 -3276 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587200 150076 587800 150078
rect -4816 150054 588740 150076
rect -4816 149818 -3694 150054
rect -3458 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587382 150054
rect 587618 149818 588740 150054
rect -4816 149734 588740 149818
rect -4816 149498 -3694 149734
rect -3458 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587382 149734
rect 587618 149498 588740 149734
rect -4816 149476 588740 149498
rect -3876 149474 -3276 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587200 149474 587800 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8576 139276 -7976 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591900 139276 592500 139278
rect -8576 139254 592500 139276
rect -8576 139018 -8394 139254
rect -8158 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 592082 139254
rect 592318 139018 592500 139254
rect -8576 138934 592500 139018
rect -8576 138698 -8394 138934
rect -8158 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 592082 138934
rect 592318 138698 592500 138934
rect -8576 138676 592500 138698
rect -8576 138674 -7976 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591900 138674 592500 138676
rect -6696 135676 -6096 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 590020 135676 590620 135678
rect -6696 135654 590620 135676
rect -6696 135418 -6514 135654
rect -6278 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590202 135654
rect 590438 135418 590620 135654
rect -6696 135334 590620 135418
rect -6696 135098 -6514 135334
rect -6278 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590202 135334
rect 590438 135098 590620 135334
rect -6696 135076 590620 135098
rect -6696 135074 -6096 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 590020 135074 590620 135076
rect -4816 132076 -4216 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588140 132076 588740 132078
rect -4816 132054 588740 132076
rect -4816 131818 -4634 132054
rect -4398 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588322 132054
rect 588558 131818 588740 132054
rect -4816 131734 588740 131818
rect -4816 131498 -4634 131734
rect -4398 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588322 131734
rect 588558 131498 588740 131734
rect -4816 131476 588740 131498
rect -4816 131474 -4216 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588140 131474 588740 131476
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -7636 121276 -7036 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590960 121276 591560 121278
rect -8576 121254 592500 121276
rect -8576 121018 -7454 121254
rect -7218 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591142 121254
rect 591378 121018 592500 121254
rect -8576 120934 592500 121018
rect -8576 120698 -7454 120934
rect -7218 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591142 120934
rect 591378 120698 592500 120934
rect -8576 120676 592500 120698
rect -7636 120674 -7036 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590960 120674 591560 120676
rect -5756 117676 -5156 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589080 117676 589680 117678
rect -6696 117654 590620 117676
rect -6696 117418 -5574 117654
rect -5338 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589262 117654
rect 589498 117418 590620 117654
rect -6696 117334 590620 117418
rect -6696 117098 -5574 117334
rect -5338 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589262 117334
rect 589498 117098 590620 117334
rect -6696 117076 590620 117098
rect -5756 117074 -5156 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589080 117074 589680 117076
rect -3876 114076 -3276 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587200 114076 587800 114078
rect -4816 114054 588740 114076
rect -4816 113818 -3694 114054
rect -3458 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587382 114054
rect 587618 113818 588740 114054
rect -4816 113734 588740 113818
rect -4816 113498 -3694 113734
rect -3458 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587382 113734
rect 587618 113498 588740 113734
rect -4816 113476 588740 113498
rect -3876 113474 -3276 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587200 113474 587800 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8576 103276 -7976 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591900 103276 592500 103278
rect -8576 103254 592500 103276
rect -8576 103018 -8394 103254
rect -8158 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 592082 103254
rect 592318 103018 592500 103254
rect -8576 102934 592500 103018
rect -8576 102698 -8394 102934
rect -8158 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 592082 102934
rect 592318 102698 592500 102934
rect -8576 102676 592500 102698
rect -8576 102674 -7976 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591900 102674 592500 102676
rect -6696 99676 -6096 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 590020 99676 590620 99678
rect -6696 99654 590620 99676
rect -6696 99418 -6514 99654
rect -6278 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590202 99654
rect 590438 99418 590620 99654
rect -6696 99334 590620 99418
rect -6696 99098 -6514 99334
rect -6278 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590202 99334
rect 590438 99098 590620 99334
rect -6696 99076 590620 99098
rect -6696 99074 -6096 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 590020 99074 590620 99076
rect -4816 96076 -4216 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588140 96076 588740 96078
rect -4816 96054 588740 96076
rect -4816 95818 -4634 96054
rect -4398 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588322 96054
rect 588558 95818 588740 96054
rect -4816 95734 588740 95818
rect -4816 95498 -4634 95734
rect -4398 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588322 95734
rect 588558 95498 588740 95734
rect -4816 95476 588740 95498
rect -4816 95474 -4216 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588140 95474 588740 95476
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -7636 85276 -7036 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590960 85276 591560 85278
rect -8576 85254 592500 85276
rect -8576 85018 -7454 85254
rect -7218 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591142 85254
rect 591378 85018 592500 85254
rect -8576 84934 592500 85018
rect -8576 84698 -7454 84934
rect -7218 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591142 84934
rect 591378 84698 592500 84934
rect -8576 84676 592500 84698
rect -7636 84674 -7036 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590960 84674 591560 84676
rect -5756 81676 -5156 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589080 81676 589680 81678
rect -6696 81654 590620 81676
rect -6696 81418 -5574 81654
rect -5338 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589262 81654
rect 589498 81418 590620 81654
rect -6696 81334 590620 81418
rect -6696 81098 -5574 81334
rect -5338 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589262 81334
rect 589498 81098 590620 81334
rect -6696 81076 590620 81098
rect -5756 81074 -5156 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589080 81074 589680 81076
rect -3876 78076 -3276 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587200 78076 587800 78078
rect -4816 78054 588740 78076
rect -4816 77818 -3694 78054
rect -3458 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587382 78054
rect 587618 77818 588740 78054
rect -4816 77734 588740 77818
rect -4816 77498 -3694 77734
rect -3458 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587382 77734
rect 587618 77498 588740 77734
rect -4816 77476 588740 77498
rect -3876 77474 -3276 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587200 77474 587800 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8576 67276 -7976 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591900 67276 592500 67278
rect -8576 67254 592500 67276
rect -8576 67018 -8394 67254
rect -8158 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 592082 67254
rect 592318 67018 592500 67254
rect -8576 66934 592500 67018
rect -8576 66698 -8394 66934
rect -8158 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 592082 66934
rect 592318 66698 592500 66934
rect -8576 66676 592500 66698
rect -8576 66674 -7976 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591900 66674 592500 66676
rect -6696 63676 -6096 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 590020 63676 590620 63678
rect -6696 63654 590620 63676
rect -6696 63418 -6514 63654
rect -6278 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590202 63654
rect 590438 63418 590620 63654
rect -6696 63334 590620 63418
rect -6696 63098 -6514 63334
rect -6278 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590202 63334
rect 590438 63098 590620 63334
rect -6696 63076 590620 63098
rect -6696 63074 -6096 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 590020 63074 590620 63076
rect -4816 60076 -4216 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588140 60076 588740 60078
rect -4816 60054 588740 60076
rect -4816 59818 -4634 60054
rect -4398 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588322 60054
rect 588558 59818 588740 60054
rect -4816 59734 588740 59818
rect -4816 59498 -4634 59734
rect -4398 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588322 59734
rect 588558 59498 588740 59734
rect -4816 59476 588740 59498
rect -4816 59474 -4216 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588140 59474 588740 59476
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -7636 49276 -7036 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590960 49276 591560 49278
rect -8576 49254 592500 49276
rect -8576 49018 -7454 49254
rect -7218 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591142 49254
rect 591378 49018 592500 49254
rect -8576 48934 592500 49018
rect -8576 48698 -7454 48934
rect -7218 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591142 48934
rect 591378 48698 592500 48934
rect -8576 48676 592500 48698
rect -7636 48674 -7036 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590960 48674 591560 48676
rect -5756 45676 -5156 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589080 45676 589680 45678
rect -6696 45654 590620 45676
rect -6696 45418 -5574 45654
rect -5338 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589262 45654
rect 589498 45418 590620 45654
rect -6696 45334 590620 45418
rect -6696 45098 -5574 45334
rect -5338 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589262 45334
rect 589498 45098 590620 45334
rect -6696 45076 590620 45098
rect -5756 45074 -5156 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589080 45074 589680 45076
rect -3876 42076 -3276 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587200 42076 587800 42078
rect -4816 42054 588740 42076
rect -4816 41818 -3694 42054
rect -3458 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587382 42054
rect 587618 41818 588740 42054
rect -4816 41734 588740 41818
rect -4816 41498 -3694 41734
rect -3458 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587382 41734
rect 587618 41498 588740 41734
rect -4816 41476 588740 41498
rect -3876 41474 -3276 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587200 41474 587800 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8576 31276 -7976 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591900 31276 592500 31278
rect -8576 31254 592500 31276
rect -8576 31018 -8394 31254
rect -8158 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 592082 31254
rect 592318 31018 592500 31254
rect -8576 30934 592500 31018
rect -8576 30698 -8394 30934
rect -8158 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 592082 30934
rect 592318 30698 592500 30934
rect -8576 30676 592500 30698
rect -8576 30674 -7976 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591900 30674 592500 30676
rect -6696 27676 -6096 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 590020 27676 590620 27678
rect -6696 27654 590620 27676
rect -6696 27418 -6514 27654
rect -6278 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590202 27654
rect 590438 27418 590620 27654
rect -6696 27334 590620 27418
rect -6696 27098 -6514 27334
rect -6278 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590202 27334
rect 590438 27098 590620 27334
rect -6696 27076 590620 27098
rect -6696 27074 -6096 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 590020 27074 590620 27076
rect -4816 24076 -4216 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588140 24076 588740 24078
rect -4816 24054 588740 24076
rect -4816 23818 -4634 24054
rect -4398 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588322 24054
rect 588558 23818 588740 24054
rect -4816 23734 588740 23818
rect -4816 23498 -4634 23734
rect -4398 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588322 23734
rect 588558 23498 588740 23734
rect -4816 23476 588740 23498
rect -4816 23474 -4216 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588140 23474 588740 23476
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -7636 13276 -7036 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590960 13276 591560 13278
rect -8576 13254 592500 13276
rect -8576 13018 -7454 13254
rect -7218 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591142 13254
rect 591378 13018 592500 13254
rect -8576 12934 592500 13018
rect -8576 12698 -7454 12934
rect -7218 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591142 12934
rect 591378 12698 592500 12934
rect -8576 12676 592500 12698
rect -7636 12674 -7036 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590960 12674 591560 12676
rect -5756 9676 -5156 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589080 9676 589680 9678
rect -6696 9654 590620 9676
rect -6696 9418 -5574 9654
rect -5338 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589262 9654
rect 589498 9418 590620 9654
rect -6696 9334 590620 9418
rect -6696 9098 -5574 9334
rect -5338 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589262 9334
rect 589498 9098 590620 9334
rect -6696 9076 590620 9098
rect -5756 9074 -5156 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589080 9074 589680 9076
rect -3876 6076 -3276 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587200 6076 587800 6078
rect -4816 6054 588740 6076
rect -4816 5818 -3694 6054
rect -3458 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587382 6054
rect 587618 5818 588740 6054
rect -4816 5734 588740 5818
rect -4816 5498 -3694 5734
rect -3458 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587382 5734
rect 587618 5498 588740 5734
rect -4816 5476 588740 5498
rect -3876 5474 -3276 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587200 5474 587800 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 4586 -2226
rect 4822 -2462 40586 -2226
rect 40822 -2462 76586 -2226
rect 76822 -2462 112586 -2226
rect 112822 -2462 148586 -2226
rect 148822 -2462 184586 -2226
rect 184822 -2462 220586 -2226
rect 220822 -2462 256586 -2226
rect 256822 -2462 292586 -2226
rect 292822 -2462 328586 -2226
rect 328822 -2462 364586 -2226
rect 364822 -2462 400586 -2226
rect 400822 -2462 436586 -2226
rect 436822 -2462 472586 -2226
rect 472822 -2462 508586 -2226
rect 508822 -2462 544586 -2226
rect 544822 -2462 580586 -2226
rect 580822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 4586 -2546
rect 4822 -2782 40586 -2546
rect 40822 -2782 76586 -2546
rect 76822 -2782 112586 -2546
rect 112822 -2782 148586 -2546
rect 148822 -2782 184586 -2546
rect 184822 -2782 220586 -2546
rect 220822 -2782 256586 -2546
rect 256822 -2782 292586 -2546
rect 292822 -2782 328586 -2546
rect 328822 -2782 364586 -2546
rect 364822 -2782 400586 -2546
rect 400822 -2782 436586 -2546
rect 436822 -2782 472586 -2546
rect 472822 -2782 508586 -2546
rect 508822 -2782 544586 -2546
rect 544822 -2782 580586 -2546
rect 580822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 22586 -3166
rect 22822 -3402 58586 -3166
rect 58822 -3402 94586 -3166
rect 94822 -3402 130586 -3166
rect 130822 -3402 166586 -3166
rect 166822 -3402 202586 -3166
rect 202822 -3402 238586 -3166
rect 238822 -3402 274586 -3166
rect 274822 -3402 310586 -3166
rect 310822 -3402 346586 -3166
rect 346822 -3402 382586 -3166
rect 382822 -3402 418586 -3166
rect 418822 -3402 454586 -3166
rect 454822 -3402 490586 -3166
rect 490822 -3402 526586 -3166
rect 526822 -3402 562586 -3166
rect 562822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 22586 -3486
rect 22822 -3722 58586 -3486
rect 58822 -3722 94586 -3486
rect 94822 -3722 130586 -3486
rect 130822 -3722 166586 -3486
rect 166822 -3722 202586 -3486
rect 202822 -3722 238586 -3486
rect 238822 -3722 274586 -3486
rect 274822 -3722 310586 -3486
rect 310822 -3722 346586 -3486
rect 346822 -3722 382586 -3486
rect 382822 -3722 418586 -3486
rect 418822 -3722 454586 -3486
rect 454822 -3722 490586 -3486
rect 490822 -3722 526586 -3486
rect 526822 -3722 562586 -3486
rect 562822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 8186 -4106
rect 8422 -4342 44186 -4106
rect 44422 -4342 80186 -4106
rect 80422 -4342 116186 -4106
rect 116422 -4342 152186 -4106
rect 152422 -4342 188186 -4106
rect 188422 -4342 224186 -4106
rect 224422 -4342 260186 -4106
rect 260422 -4342 296186 -4106
rect 296422 -4342 332186 -4106
rect 332422 -4342 368186 -4106
rect 368422 -4342 404186 -4106
rect 404422 -4342 440186 -4106
rect 440422 -4342 476186 -4106
rect 476422 -4342 512186 -4106
rect 512422 -4342 548186 -4106
rect 548422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 8186 -4426
rect 8422 -4662 44186 -4426
rect 44422 -4662 80186 -4426
rect 80422 -4662 116186 -4426
rect 116422 -4662 152186 -4426
rect 152422 -4662 188186 -4426
rect 188422 -4662 224186 -4426
rect 224422 -4662 260186 -4426
rect 260422 -4662 296186 -4426
rect 296422 -4662 332186 -4426
rect 332422 -4662 368186 -4426
rect 368422 -4662 404186 -4426
rect 404422 -4662 440186 -4426
rect 440422 -4662 476186 -4426
rect 476422 -4662 512186 -4426
rect 512422 -4662 548186 -4426
rect 548422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 26186 -5046
rect 26422 -5282 62186 -5046
rect 62422 -5282 98186 -5046
rect 98422 -5282 134186 -5046
rect 134422 -5282 170186 -5046
rect 170422 -5282 206186 -5046
rect 206422 -5282 242186 -5046
rect 242422 -5282 278186 -5046
rect 278422 -5282 314186 -5046
rect 314422 -5282 350186 -5046
rect 350422 -5282 386186 -5046
rect 386422 -5282 422186 -5046
rect 422422 -5282 458186 -5046
rect 458422 -5282 494186 -5046
rect 494422 -5282 530186 -5046
rect 530422 -5282 566186 -5046
rect 566422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 26186 -5366
rect 26422 -5602 62186 -5366
rect 62422 -5602 98186 -5366
rect 98422 -5602 134186 -5366
rect 134422 -5602 170186 -5366
rect 170422 -5602 206186 -5366
rect 206422 -5602 242186 -5366
rect 242422 -5602 278186 -5366
rect 278422 -5602 314186 -5366
rect 314422 -5602 350186 -5366
rect 350422 -5602 386186 -5366
rect 386422 -5602 422186 -5366
rect 422422 -5602 458186 -5366
rect 458422 -5602 494186 -5366
rect 494422 -5602 530186 -5366
rect 530422 -5602 566186 -5366
rect 566422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 11786 -5986
rect 12022 -6222 47786 -5986
rect 48022 -6222 83786 -5986
rect 84022 -6222 119786 -5986
rect 120022 -6222 155786 -5986
rect 156022 -6222 191786 -5986
rect 192022 -6222 227786 -5986
rect 228022 -6222 263786 -5986
rect 264022 -6222 299786 -5986
rect 300022 -6222 335786 -5986
rect 336022 -6222 371786 -5986
rect 372022 -6222 407786 -5986
rect 408022 -6222 443786 -5986
rect 444022 -6222 479786 -5986
rect 480022 -6222 515786 -5986
rect 516022 -6222 551786 -5986
rect 552022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 11786 -6306
rect 12022 -6542 47786 -6306
rect 48022 -6542 83786 -6306
rect 84022 -6542 119786 -6306
rect 120022 -6542 155786 -6306
rect 156022 -6542 191786 -6306
rect 192022 -6542 227786 -6306
rect 228022 -6542 263786 -6306
rect 264022 -6542 299786 -6306
rect 300022 -6542 335786 -6306
rect 336022 -6542 371786 -6306
rect 372022 -6542 407786 -6306
rect 408022 -6542 443786 -6306
rect 444022 -6542 479786 -6306
rect 480022 -6542 515786 -6306
rect 516022 -6542 551786 -6306
rect 552022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 29786 -6926
rect 30022 -7162 65786 -6926
rect 66022 -7162 101786 -6926
rect 102022 -7162 137786 -6926
rect 138022 -7162 173786 -6926
rect 174022 -7162 209786 -6926
rect 210022 -7162 245786 -6926
rect 246022 -7162 281786 -6926
rect 282022 -7162 317786 -6926
rect 318022 -7162 353786 -6926
rect 354022 -7162 389786 -6926
rect 390022 -7162 425786 -6926
rect 426022 -7162 461786 -6926
rect 462022 -7162 497786 -6926
rect 498022 -7162 533786 -6926
rect 534022 -7162 569786 -6926
rect 570022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 29786 -7246
rect 30022 -7482 65786 -7246
rect 66022 -7482 101786 -7246
rect 102022 -7482 137786 -7246
rect 138022 -7482 173786 -7246
rect 174022 -7482 209786 -7246
rect 210022 -7482 245786 -7246
rect 246022 -7482 281786 -7246
rect 282022 -7482 317786 -7246
rect 318022 -7482 353786 -7246
rect 354022 -7482 389786 -7246
rect 390022 -7482 425786 -7246
rect 426022 -7482 461786 -7246
rect 462022 -7482 497786 -7246
rect 498022 -7482 533786 -7246
rect 534022 -7482 569786 -7246
rect 570022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
use accelerator_top  mprj
timestamp 1608101209
transform 1 0 155000 0 1 175000
box 0 0 234658 236802
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1608252747
<< obsli1 >>
rect 1104 2159 289064 289969
<< obsm1 >>
rect 842 1028 289418 290000
<< metal2 >>
rect 5354 291595 5410 292395
rect 16026 291595 16082 292395
rect 26790 291595 26846 292395
rect 37554 291595 37610 292395
rect 48318 291595 48374 292395
rect 59082 291595 59138 292395
rect 69846 291595 69902 292395
rect 80518 291595 80574 292395
rect 91282 291595 91338 292395
rect 102046 291595 102102 292395
rect 112810 291595 112866 292395
rect 123574 291595 123630 292395
rect 134338 291595 134394 292395
rect 145102 291595 145158 292395
rect 155774 291595 155830 292395
rect 166538 291595 166594 292395
rect 177302 291595 177358 292395
rect 188066 291595 188122 292395
rect 198830 291595 198886 292395
rect 209594 291595 209650 292395
rect 220358 291595 220414 292395
rect 231030 291595 231086 292395
rect 241794 291595 241850 292395
rect 252558 291595 252614 292395
rect 263322 291595 263378 292395
rect 274086 291595 274142 292395
rect 284850 291595 284906 292395
rect 294 0 350 800
rect 846 0 902 800
rect 1398 0 1454 800
rect 2042 0 2098 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3790 0 3846 800
rect 4434 0 4490 800
rect 4986 0 5042 800
rect 5538 0 5594 800
rect 6182 0 6238 800
rect 6734 0 6790 800
rect 7378 0 7434 800
rect 7930 0 7986 800
rect 8574 0 8630 800
rect 9126 0 9182 800
rect 9770 0 9826 800
rect 10322 0 10378 800
rect 10874 0 10930 800
rect 11518 0 11574 800
rect 12070 0 12126 800
rect 12714 0 12770 800
rect 13266 0 13322 800
rect 13910 0 13966 800
rect 14462 0 14518 800
rect 15014 0 15070 800
rect 15658 0 15714 800
rect 16210 0 16266 800
rect 16854 0 16910 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18602 0 18658 800
rect 19246 0 19302 800
rect 19798 0 19854 800
rect 20350 0 20406 800
rect 20994 0 21050 800
rect 21546 0 21602 800
rect 22190 0 22246 800
rect 22742 0 22798 800
rect 23386 0 23442 800
rect 23938 0 23994 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25686 0 25742 800
rect 26330 0 26386 800
rect 26882 0 26938 800
rect 27526 0 27582 800
rect 28078 0 28134 800
rect 28722 0 28778 800
rect 29274 0 29330 800
rect 29826 0 29882 800
rect 30470 0 30526 800
rect 31022 0 31078 800
rect 31666 0 31722 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33414 0 33470 800
rect 34058 0 34114 800
rect 34610 0 34666 800
rect 35162 0 35218 800
rect 35806 0 35862 800
rect 36358 0 36414 800
rect 37002 0 37058 800
rect 37554 0 37610 800
rect 38198 0 38254 800
rect 38750 0 38806 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40498 0 40554 800
rect 41142 0 41198 800
rect 41694 0 41750 800
rect 42338 0 42394 800
rect 42890 0 42946 800
rect 43534 0 43590 800
rect 44086 0 44142 800
rect 44638 0 44694 800
rect 45282 0 45338 800
rect 45834 0 45890 800
rect 46478 0 46534 800
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 48226 0 48282 800
rect 48778 0 48834 800
rect 49422 0 49478 800
rect 49974 0 50030 800
rect 50618 0 50674 800
rect 51170 0 51226 800
rect 51814 0 51870 800
rect 52366 0 52422 800
rect 53010 0 53066 800
rect 53562 0 53618 800
rect 54114 0 54170 800
rect 54758 0 54814 800
rect 55310 0 55366 800
rect 55954 0 56010 800
rect 56506 0 56562 800
rect 57150 0 57206 800
rect 57702 0 57758 800
rect 58346 0 58402 800
rect 58898 0 58954 800
rect 59450 0 59506 800
rect 60094 0 60150 800
rect 60646 0 60702 800
rect 61290 0 61346 800
rect 61842 0 61898 800
rect 62486 0 62542 800
rect 63038 0 63094 800
rect 63590 0 63646 800
rect 64234 0 64290 800
rect 64786 0 64842 800
rect 65430 0 65486 800
rect 65982 0 66038 800
rect 66626 0 66682 800
rect 67178 0 67234 800
rect 67822 0 67878 800
rect 68374 0 68430 800
rect 68926 0 68982 800
rect 69570 0 69626 800
rect 70122 0 70178 800
rect 70766 0 70822 800
rect 71318 0 71374 800
rect 71962 0 72018 800
rect 72514 0 72570 800
rect 73066 0 73122 800
rect 73710 0 73766 800
rect 74262 0 74318 800
rect 74906 0 74962 800
rect 75458 0 75514 800
rect 76102 0 76158 800
rect 76654 0 76710 800
rect 77298 0 77354 800
rect 77850 0 77906 800
rect 78402 0 78458 800
rect 79046 0 79102 800
rect 79598 0 79654 800
rect 80242 0 80298 800
rect 80794 0 80850 800
rect 81438 0 81494 800
rect 81990 0 82046 800
rect 82542 0 82598 800
rect 83186 0 83242 800
rect 83738 0 83794 800
rect 84382 0 84438 800
rect 84934 0 84990 800
rect 85578 0 85634 800
rect 86130 0 86186 800
rect 86774 0 86830 800
rect 87326 0 87382 800
rect 87878 0 87934 800
rect 88522 0 88578 800
rect 89074 0 89130 800
rect 89718 0 89774 800
rect 90270 0 90326 800
rect 90914 0 90970 800
rect 91466 0 91522 800
rect 92110 0 92166 800
rect 92662 0 92718 800
rect 93214 0 93270 800
rect 93858 0 93914 800
rect 94410 0 94466 800
rect 95054 0 95110 800
rect 95606 0 95662 800
rect 96250 0 96306 800
rect 96802 0 96858 800
rect 97354 0 97410 800
rect 97998 0 98054 800
rect 98550 0 98606 800
rect 99194 0 99250 800
rect 99746 0 99802 800
rect 100390 0 100446 800
rect 100942 0 100998 800
rect 101586 0 101642 800
rect 102138 0 102194 800
rect 102690 0 102746 800
rect 103334 0 103390 800
rect 103886 0 103942 800
rect 104530 0 104586 800
rect 105082 0 105138 800
rect 105726 0 105782 800
rect 106278 0 106334 800
rect 106830 0 106886 800
rect 107474 0 107530 800
rect 108026 0 108082 800
rect 108670 0 108726 800
rect 109222 0 109278 800
rect 109866 0 109922 800
rect 110418 0 110474 800
rect 111062 0 111118 800
rect 111614 0 111670 800
rect 112166 0 112222 800
rect 112810 0 112866 800
rect 113362 0 113418 800
rect 114006 0 114062 800
rect 114558 0 114614 800
rect 115202 0 115258 800
rect 115754 0 115810 800
rect 116398 0 116454 800
rect 116950 0 117006 800
rect 117502 0 117558 800
rect 118146 0 118202 800
rect 118698 0 118754 800
rect 119342 0 119398 800
rect 119894 0 119950 800
rect 120538 0 120594 800
rect 121090 0 121146 800
rect 121642 0 121698 800
rect 122286 0 122342 800
rect 122838 0 122894 800
rect 123482 0 123538 800
rect 124034 0 124090 800
rect 124678 0 124734 800
rect 125230 0 125286 800
rect 125874 0 125930 800
rect 126426 0 126482 800
rect 126978 0 127034 800
rect 127622 0 127678 800
rect 128174 0 128230 800
rect 128818 0 128874 800
rect 129370 0 129426 800
rect 130014 0 130070 800
rect 130566 0 130622 800
rect 131118 0 131174 800
rect 131762 0 131818 800
rect 132314 0 132370 800
rect 132958 0 133014 800
rect 133510 0 133566 800
rect 134154 0 134210 800
rect 134706 0 134762 800
rect 135350 0 135406 800
rect 135902 0 135958 800
rect 136454 0 136510 800
rect 137098 0 137154 800
rect 137650 0 137706 800
rect 138294 0 138350 800
rect 138846 0 138902 800
rect 139490 0 139546 800
rect 140042 0 140098 800
rect 140594 0 140650 800
rect 141238 0 141294 800
rect 141790 0 141846 800
rect 142434 0 142490 800
rect 142986 0 143042 800
rect 143630 0 143686 800
rect 144182 0 144238 800
rect 144826 0 144882 800
rect 145378 0 145434 800
rect 145930 0 145986 800
rect 146574 0 146630 800
rect 147126 0 147182 800
rect 147770 0 147826 800
rect 148322 0 148378 800
rect 148966 0 149022 800
rect 149518 0 149574 800
rect 150162 0 150218 800
rect 150714 0 150770 800
rect 151266 0 151322 800
rect 151910 0 151966 800
rect 152462 0 152518 800
rect 153106 0 153162 800
rect 153658 0 153714 800
rect 154302 0 154358 800
rect 154854 0 154910 800
rect 155406 0 155462 800
rect 156050 0 156106 800
rect 156602 0 156658 800
rect 157246 0 157302 800
rect 157798 0 157854 800
rect 158442 0 158498 800
rect 158994 0 159050 800
rect 159638 0 159694 800
rect 160190 0 160246 800
rect 160742 0 160798 800
rect 161386 0 161442 800
rect 161938 0 161994 800
rect 162582 0 162638 800
rect 163134 0 163190 800
rect 163778 0 163834 800
rect 164330 0 164386 800
rect 164882 0 164938 800
rect 165526 0 165582 800
rect 166078 0 166134 800
rect 166722 0 166778 800
rect 167274 0 167330 800
rect 167918 0 167974 800
rect 168470 0 168526 800
rect 169114 0 169170 800
rect 169666 0 169722 800
rect 170218 0 170274 800
rect 170862 0 170918 800
rect 171414 0 171470 800
rect 172058 0 172114 800
rect 172610 0 172666 800
rect 173254 0 173310 800
rect 173806 0 173862 800
rect 174450 0 174506 800
rect 175002 0 175058 800
rect 175554 0 175610 800
rect 176198 0 176254 800
rect 176750 0 176806 800
rect 177394 0 177450 800
rect 177946 0 178002 800
rect 178590 0 178646 800
rect 179142 0 179198 800
rect 179694 0 179750 800
rect 180338 0 180394 800
rect 180890 0 180946 800
rect 181534 0 181590 800
rect 182086 0 182142 800
rect 182730 0 182786 800
rect 183282 0 183338 800
rect 183926 0 183982 800
rect 184478 0 184534 800
rect 185030 0 185086 800
rect 185674 0 185730 800
rect 186226 0 186282 800
rect 186870 0 186926 800
rect 187422 0 187478 800
rect 188066 0 188122 800
rect 188618 0 188674 800
rect 189170 0 189226 800
rect 189814 0 189870 800
rect 190366 0 190422 800
rect 191010 0 191066 800
rect 191562 0 191618 800
rect 192206 0 192262 800
rect 192758 0 192814 800
rect 193402 0 193458 800
rect 193954 0 194010 800
rect 194506 0 194562 800
rect 195150 0 195206 800
rect 195702 0 195758 800
rect 196346 0 196402 800
rect 196898 0 196954 800
rect 197542 0 197598 800
rect 198094 0 198150 800
rect 198646 0 198702 800
rect 199290 0 199346 800
rect 199842 0 199898 800
rect 200486 0 200542 800
rect 201038 0 201094 800
rect 201682 0 201738 800
rect 202234 0 202290 800
rect 202878 0 202934 800
rect 203430 0 203486 800
rect 203982 0 204038 800
rect 204626 0 204682 800
rect 205178 0 205234 800
rect 205822 0 205878 800
rect 206374 0 206430 800
rect 207018 0 207074 800
rect 207570 0 207626 800
rect 208214 0 208270 800
rect 208766 0 208822 800
rect 209318 0 209374 800
rect 209962 0 210018 800
rect 210514 0 210570 800
rect 211158 0 211214 800
rect 211710 0 211766 800
rect 212354 0 212410 800
rect 212906 0 212962 800
rect 213458 0 213514 800
rect 214102 0 214158 800
rect 214654 0 214710 800
rect 215298 0 215354 800
rect 215850 0 215906 800
rect 216494 0 216550 800
rect 217046 0 217102 800
rect 217690 0 217746 800
rect 218242 0 218298 800
rect 218794 0 218850 800
rect 219438 0 219494 800
rect 219990 0 220046 800
rect 220634 0 220690 800
rect 221186 0 221242 800
rect 221830 0 221886 800
rect 222382 0 222438 800
rect 222934 0 222990 800
rect 223578 0 223634 800
rect 224130 0 224186 800
rect 224774 0 224830 800
rect 225326 0 225382 800
rect 225970 0 226026 800
rect 226522 0 226578 800
rect 227166 0 227222 800
rect 227718 0 227774 800
rect 228270 0 228326 800
rect 228914 0 228970 800
rect 229466 0 229522 800
rect 230110 0 230166 800
rect 230662 0 230718 800
rect 231306 0 231362 800
rect 231858 0 231914 800
rect 232502 0 232558 800
rect 233054 0 233110 800
rect 233606 0 233662 800
rect 234250 0 234306 800
rect 234802 0 234858 800
rect 235446 0 235502 800
rect 235998 0 236054 800
rect 236642 0 236698 800
rect 237194 0 237250 800
rect 237746 0 237802 800
rect 238390 0 238446 800
rect 238942 0 238998 800
rect 239586 0 239642 800
rect 240138 0 240194 800
rect 240782 0 240838 800
rect 241334 0 241390 800
rect 241978 0 242034 800
rect 242530 0 242586 800
rect 243082 0 243138 800
rect 243726 0 243782 800
rect 244278 0 244334 800
rect 244922 0 244978 800
rect 245474 0 245530 800
rect 246118 0 246174 800
rect 246670 0 246726 800
rect 247222 0 247278 800
rect 247866 0 247922 800
rect 248418 0 248474 800
rect 249062 0 249118 800
rect 249614 0 249670 800
rect 250258 0 250314 800
rect 250810 0 250866 800
rect 251454 0 251510 800
rect 252006 0 252062 800
rect 252558 0 252614 800
rect 253202 0 253258 800
rect 253754 0 253810 800
rect 254398 0 254454 800
rect 254950 0 255006 800
rect 255594 0 255650 800
rect 256146 0 256202 800
rect 256698 0 256754 800
rect 257342 0 257398 800
rect 257894 0 257950 800
rect 258538 0 258594 800
rect 259090 0 259146 800
rect 259734 0 259790 800
rect 260286 0 260342 800
rect 260930 0 260986 800
rect 261482 0 261538 800
rect 262034 0 262090 800
rect 262678 0 262734 800
rect 263230 0 263286 800
rect 263874 0 263930 800
rect 264426 0 264482 800
rect 265070 0 265126 800
rect 265622 0 265678 800
rect 266266 0 266322 800
rect 266818 0 266874 800
rect 267370 0 267426 800
rect 268014 0 268070 800
rect 268566 0 268622 800
rect 269210 0 269266 800
rect 269762 0 269818 800
rect 270406 0 270462 800
rect 270958 0 271014 800
rect 271510 0 271566 800
rect 272154 0 272210 800
rect 272706 0 272762 800
rect 273350 0 273406 800
rect 273902 0 273958 800
rect 274546 0 274602 800
rect 275098 0 275154 800
rect 275742 0 275798 800
rect 276294 0 276350 800
rect 276846 0 276902 800
rect 277490 0 277546 800
rect 278042 0 278098 800
rect 278686 0 278742 800
rect 279238 0 279294 800
rect 279882 0 279938 800
rect 280434 0 280490 800
rect 280986 0 281042 800
rect 281630 0 281686 800
rect 282182 0 282238 800
rect 282826 0 282882 800
rect 283378 0 283434 800
rect 284022 0 284078 800
rect 284574 0 284630 800
rect 285218 0 285274 800
rect 285770 0 285826 800
rect 286322 0 286378 800
rect 286966 0 287022 800
rect 287518 0 287574 800
rect 288162 0 288218 800
rect 288714 0 288770 800
rect 289358 0 289414 800
rect 289910 0 289966 800
<< obsm2 >>
rect 294 291539 5298 291595
rect 5466 291539 15970 291595
rect 16138 291539 26734 291595
rect 26902 291539 37498 291595
rect 37666 291539 48262 291595
rect 48430 291539 59026 291595
rect 59194 291539 69790 291595
rect 69958 291539 80462 291595
rect 80630 291539 91226 291595
rect 91394 291539 101990 291595
rect 102158 291539 112754 291595
rect 112922 291539 123518 291595
rect 123686 291539 134282 291595
rect 134450 291539 145046 291595
rect 145214 291539 155718 291595
rect 155886 291539 166482 291595
rect 166650 291539 177246 291595
rect 177414 291539 188010 291595
rect 188178 291539 198774 291595
rect 198942 291539 209538 291595
rect 209706 291539 220302 291595
rect 220470 291539 230974 291595
rect 231142 291539 241738 291595
rect 241906 291539 252502 291595
rect 252670 291539 263266 291595
rect 263434 291539 274030 291595
rect 274198 291539 284794 291595
rect 284962 291539 289412 291595
rect 294 856 289412 291539
rect 406 800 790 856
rect 958 800 1342 856
rect 1510 800 1986 856
rect 2154 800 2538 856
rect 2706 800 3182 856
rect 3350 800 3734 856
rect 3902 800 4378 856
rect 4546 800 4930 856
rect 5098 800 5482 856
rect 5650 800 6126 856
rect 6294 800 6678 856
rect 6846 800 7322 856
rect 7490 800 7874 856
rect 8042 800 8518 856
rect 8686 800 9070 856
rect 9238 800 9714 856
rect 9882 800 10266 856
rect 10434 800 10818 856
rect 10986 800 11462 856
rect 11630 800 12014 856
rect 12182 800 12658 856
rect 12826 800 13210 856
rect 13378 800 13854 856
rect 14022 800 14406 856
rect 14574 800 14958 856
rect 15126 800 15602 856
rect 15770 800 16154 856
rect 16322 800 16798 856
rect 16966 800 17350 856
rect 17518 800 17994 856
rect 18162 800 18546 856
rect 18714 800 19190 856
rect 19358 800 19742 856
rect 19910 800 20294 856
rect 20462 800 20938 856
rect 21106 800 21490 856
rect 21658 800 22134 856
rect 22302 800 22686 856
rect 22854 800 23330 856
rect 23498 800 23882 856
rect 24050 800 24434 856
rect 24602 800 25078 856
rect 25246 800 25630 856
rect 25798 800 26274 856
rect 26442 800 26826 856
rect 26994 800 27470 856
rect 27638 800 28022 856
rect 28190 800 28666 856
rect 28834 800 29218 856
rect 29386 800 29770 856
rect 29938 800 30414 856
rect 30582 800 30966 856
rect 31134 800 31610 856
rect 31778 800 32162 856
rect 32330 800 32806 856
rect 32974 800 33358 856
rect 33526 800 34002 856
rect 34170 800 34554 856
rect 34722 800 35106 856
rect 35274 800 35750 856
rect 35918 800 36302 856
rect 36470 800 36946 856
rect 37114 800 37498 856
rect 37666 800 38142 856
rect 38310 800 38694 856
rect 38862 800 39246 856
rect 39414 800 39890 856
rect 40058 800 40442 856
rect 40610 800 41086 856
rect 41254 800 41638 856
rect 41806 800 42282 856
rect 42450 800 42834 856
rect 43002 800 43478 856
rect 43646 800 44030 856
rect 44198 800 44582 856
rect 44750 800 45226 856
rect 45394 800 45778 856
rect 45946 800 46422 856
rect 46590 800 46974 856
rect 47142 800 47618 856
rect 47786 800 48170 856
rect 48338 800 48722 856
rect 48890 800 49366 856
rect 49534 800 49918 856
rect 50086 800 50562 856
rect 50730 800 51114 856
rect 51282 800 51758 856
rect 51926 800 52310 856
rect 52478 800 52954 856
rect 53122 800 53506 856
rect 53674 800 54058 856
rect 54226 800 54702 856
rect 54870 800 55254 856
rect 55422 800 55898 856
rect 56066 800 56450 856
rect 56618 800 57094 856
rect 57262 800 57646 856
rect 57814 800 58290 856
rect 58458 800 58842 856
rect 59010 800 59394 856
rect 59562 800 60038 856
rect 60206 800 60590 856
rect 60758 800 61234 856
rect 61402 800 61786 856
rect 61954 800 62430 856
rect 62598 800 62982 856
rect 63150 800 63534 856
rect 63702 800 64178 856
rect 64346 800 64730 856
rect 64898 800 65374 856
rect 65542 800 65926 856
rect 66094 800 66570 856
rect 66738 800 67122 856
rect 67290 800 67766 856
rect 67934 800 68318 856
rect 68486 800 68870 856
rect 69038 800 69514 856
rect 69682 800 70066 856
rect 70234 800 70710 856
rect 70878 800 71262 856
rect 71430 800 71906 856
rect 72074 800 72458 856
rect 72626 800 73010 856
rect 73178 800 73654 856
rect 73822 800 74206 856
rect 74374 800 74850 856
rect 75018 800 75402 856
rect 75570 800 76046 856
rect 76214 800 76598 856
rect 76766 800 77242 856
rect 77410 800 77794 856
rect 77962 800 78346 856
rect 78514 800 78990 856
rect 79158 800 79542 856
rect 79710 800 80186 856
rect 80354 800 80738 856
rect 80906 800 81382 856
rect 81550 800 81934 856
rect 82102 800 82486 856
rect 82654 800 83130 856
rect 83298 800 83682 856
rect 83850 800 84326 856
rect 84494 800 84878 856
rect 85046 800 85522 856
rect 85690 800 86074 856
rect 86242 800 86718 856
rect 86886 800 87270 856
rect 87438 800 87822 856
rect 87990 800 88466 856
rect 88634 800 89018 856
rect 89186 800 89662 856
rect 89830 800 90214 856
rect 90382 800 90858 856
rect 91026 800 91410 856
rect 91578 800 92054 856
rect 92222 800 92606 856
rect 92774 800 93158 856
rect 93326 800 93802 856
rect 93970 800 94354 856
rect 94522 800 94998 856
rect 95166 800 95550 856
rect 95718 800 96194 856
rect 96362 800 96746 856
rect 96914 800 97298 856
rect 97466 800 97942 856
rect 98110 800 98494 856
rect 98662 800 99138 856
rect 99306 800 99690 856
rect 99858 800 100334 856
rect 100502 800 100886 856
rect 101054 800 101530 856
rect 101698 800 102082 856
rect 102250 800 102634 856
rect 102802 800 103278 856
rect 103446 800 103830 856
rect 103998 800 104474 856
rect 104642 800 105026 856
rect 105194 800 105670 856
rect 105838 800 106222 856
rect 106390 800 106774 856
rect 106942 800 107418 856
rect 107586 800 107970 856
rect 108138 800 108614 856
rect 108782 800 109166 856
rect 109334 800 109810 856
rect 109978 800 110362 856
rect 110530 800 111006 856
rect 111174 800 111558 856
rect 111726 800 112110 856
rect 112278 800 112754 856
rect 112922 800 113306 856
rect 113474 800 113950 856
rect 114118 800 114502 856
rect 114670 800 115146 856
rect 115314 800 115698 856
rect 115866 800 116342 856
rect 116510 800 116894 856
rect 117062 800 117446 856
rect 117614 800 118090 856
rect 118258 800 118642 856
rect 118810 800 119286 856
rect 119454 800 119838 856
rect 120006 800 120482 856
rect 120650 800 121034 856
rect 121202 800 121586 856
rect 121754 800 122230 856
rect 122398 800 122782 856
rect 122950 800 123426 856
rect 123594 800 123978 856
rect 124146 800 124622 856
rect 124790 800 125174 856
rect 125342 800 125818 856
rect 125986 800 126370 856
rect 126538 800 126922 856
rect 127090 800 127566 856
rect 127734 800 128118 856
rect 128286 800 128762 856
rect 128930 800 129314 856
rect 129482 800 129958 856
rect 130126 800 130510 856
rect 130678 800 131062 856
rect 131230 800 131706 856
rect 131874 800 132258 856
rect 132426 800 132902 856
rect 133070 800 133454 856
rect 133622 800 134098 856
rect 134266 800 134650 856
rect 134818 800 135294 856
rect 135462 800 135846 856
rect 136014 800 136398 856
rect 136566 800 137042 856
rect 137210 800 137594 856
rect 137762 800 138238 856
rect 138406 800 138790 856
rect 138958 800 139434 856
rect 139602 800 139986 856
rect 140154 800 140538 856
rect 140706 800 141182 856
rect 141350 800 141734 856
rect 141902 800 142378 856
rect 142546 800 142930 856
rect 143098 800 143574 856
rect 143742 800 144126 856
rect 144294 800 144770 856
rect 144938 800 145322 856
rect 145490 800 145874 856
rect 146042 800 146518 856
rect 146686 800 147070 856
rect 147238 800 147714 856
rect 147882 800 148266 856
rect 148434 800 148910 856
rect 149078 800 149462 856
rect 149630 800 150106 856
rect 150274 800 150658 856
rect 150826 800 151210 856
rect 151378 800 151854 856
rect 152022 800 152406 856
rect 152574 800 153050 856
rect 153218 800 153602 856
rect 153770 800 154246 856
rect 154414 800 154798 856
rect 154966 800 155350 856
rect 155518 800 155994 856
rect 156162 800 156546 856
rect 156714 800 157190 856
rect 157358 800 157742 856
rect 157910 800 158386 856
rect 158554 800 158938 856
rect 159106 800 159582 856
rect 159750 800 160134 856
rect 160302 800 160686 856
rect 160854 800 161330 856
rect 161498 800 161882 856
rect 162050 800 162526 856
rect 162694 800 163078 856
rect 163246 800 163722 856
rect 163890 800 164274 856
rect 164442 800 164826 856
rect 164994 800 165470 856
rect 165638 800 166022 856
rect 166190 800 166666 856
rect 166834 800 167218 856
rect 167386 800 167862 856
rect 168030 800 168414 856
rect 168582 800 169058 856
rect 169226 800 169610 856
rect 169778 800 170162 856
rect 170330 800 170806 856
rect 170974 800 171358 856
rect 171526 800 172002 856
rect 172170 800 172554 856
rect 172722 800 173198 856
rect 173366 800 173750 856
rect 173918 800 174394 856
rect 174562 800 174946 856
rect 175114 800 175498 856
rect 175666 800 176142 856
rect 176310 800 176694 856
rect 176862 800 177338 856
rect 177506 800 177890 856
rect 178058 800 178534 856
rect 178702 800 179086 856
rect 179254 800 179638 856
rect 179806 800 180282 856
rect 180450 800 180834 856
rect 181002 800 181478 856
rect 181646 800 182030 856
rect 182198 800 182674 856
rect 182842 800 183226 856
rect 183394 800 183870 856
rect 184038 800 184422 856
rect 184590 800 184974 856
rect 185142 800 185618 856
rect 185786 800 186170 856
rect 186338 800 186814 856
rect 186982 800 187366 856
rect 187534 800 188010 856
rect 188178 800 188562 856
rect 188730 800 189114 856
rect 189282 800 189758 856
rect 189926 800 190310 856
rect 190478 800 190954 856
rect 191122 800 191506 856
rect 191674 800 192150 856
rect 192318 800 192702 856
rect 192870 800 193346 856
rect 193514 800 193898 856
rect 194066 800 194450 856
rect 194618 800 195094 856
rect 195262 800 195646 856
rect 195814 800 196290 856
rect 196458 800 196842 856
rect 197010 800 197486 856
rect 197654 800 198038 856
rect 198206 800 198590 856
rect 198758 800 199234 856
rect 199402 800 199786 856
rect 199954 800 200430 856
rect 200598 800 200982 856
rect 201150 800 201626 856
rect 201794 800 202178 856
rect 202346 800 202822 856
rect 202990 800 203374 856
rect 203542 800 203926 856
rect 204094 800 204570 856
rect 204738 800 205122 856
rect 205290 800 205766 856
rect 205934 800 206318 856
rect 206486 800 206962 856
rect 207130 800 207514 856
rect 207682 800 208158 856
rect 208326 800 208710 856
rect 208878 800 209262 856
rect 209430 800 209906 856
rect 210074 800 210458 856
rect 210626 800 211102 856
rect 211270 800 211654 856
rect 211822 800 212298 856
rect 212466 800 212850 856
rect 213018 800 213402 856
rect 213570 800 214046 856
rect 214214 800 214598 856
rect 214766 800 215242 856
rect 215410 800 215794 856
rect 215962 800 216438 856
rect 216606 800 216990 856
rect 217158 800 217634 856
rect 217802 800 218186 856
rect 218354 800 218738 856
rect 218906 800 219382 856
rect 219550 800 219934 856
rect 220102 800 220578 856
rect 220746 800 221130 856
rect 221298 800 221774 856
rect 221942 800 222326 856
rect 222494 800 222878 856
rect 223046 800 223522 856
rect 223690 800 224074 856
rect 224242 800 224718 856
rect 224886 800 225270 856
rect 225438 800 225914 856
rect 226082 800 226466 856
rect 226634 800 227110 856
rect 227278 800 227662 856
rect 227830 800 228214 856
rect 228382 800 228858 856
rect 229026 800 229410 856
rect 229578 800 230054 856
rect 230222 800 230606 856
rect 230774 800 231250 856
rect 231418 800 231802 856
rect 231970 800 232446 856
rect 232614 800 232998 856
rect 233166 800 233550 856
rect 233718 800 234194 856
rect 234362 800 234746 856
rect 234914 800 235390 856
rect 235558 800 235942 856
rect 236110 800 236586 856
rect 236754 800 237138 856
rect 237306 800 237690 856
rect 237858 800 238334 856
rect 238502 800 238886 856
rect 239054 800 239530 856
rect 239698 800 240082 856
rect 240250 800 240726 856
rect 240894 800 241278 856
rect 241446 800 241922 856
rect 242090 800 242474 856
rect 242642 800 243026 856
rect 243194 800 243670 856
rect 243838 800 244222 856
rect 244390 800 244866 856
rect 245034 800 245418 856
rect 245586 800 246062 856
rect 246230 800 246614 856
rect 246782 800 247166 856
rect 247334 800 247810 856
rect 247978 800 248362 856
rect 248530 800 249006 856
rect 249174 800 249558 856
rect 249726 800 250202 856
rect 250370 800 250754 856
rect 250922 800 251398 856
rect 251566 800 251950 856
rect 252118 800 252502 856
rect 252670 800 253146 856
rect 253314 800 253698 856
rect 253866 800 254342 856
rect 254510 800 254894 856
rect 255062 800 255538 856
rect 255706 800 256090 856
rect 256258 800 256642 856
rect 256810 800 257286 856
rect 257454 800 257838 856
rect 258006 800 258482 856
rect 258650 800 259034 856
rect 259202 800 259678 856
rect 259846 800 260230 856
rect 260398 800 260874 856
rect 261042 800 261426 856
rect 261594 800 261978 856
rect 262146 800 262622 856
rect 262790 800 263174 856
rect 263342 800 263818 856
rect 263986 800 264370 856
rect 264538 800 265014 856
rect 265182 800 265566 856
rect 265734 800 266210 856
rect 266378 800 266762 856
rect 266930 800 267314 856
rect 267482 800 267958 856
rect 268126 800 268510 856
rect 268678 800 269154 856
rect 269322 800 269706 856
rect 269874 800 270350 856
rect 270518 800 270902 856
rect 271070 800 271454 856
rect 271622 800 272098 856
rect 272266 800 272650 856
rect 272818 800 273294 856
rect 273462 800 273846 856
rect 274014 800 274490 856
rect 274658 800 275042 856
rect 275210 800 275686 856
rect 275854 800 276238 856
rect 276406 800 276790 856
rect 276958 800 277434 856
rect 277602 800 277986 856
rect 278154 800 278630 856
rect 278798 800 279182 856
rect 279350 800 279826 856
rect 279994 800 280378 856
rect 280546 800 280930 856
rect 281098 800 281574 856
rect 281742 800 282126 856
rect 282294 800 282770 856
rect 282938 800 283322 856
rect 283490 800 283966 856
rect 284134 800 284518 856
rect 284686 800 285162 856
rect 285330 800 285714 856
rect 285882 800 286266 856
rect 286434 800 286910 856
rect 287078 800 287462 856
rect 287630 800 288106 856
rect 288274 800 288658 856
rect 288826 800 289302 856
<< metal3 >>
rect 289451 289008 290251 289128
rect 0 288736 800 288856
rect 289451 282480 290251 282600
rect 0 281800 800 281920
rect 289451 275952 290251 276072
rect 0 274864 800 274984
rect 289451 269424 290251 269544
rect 0 267928 800 268048
rect 289451 263032 290251 263152
rect 0 260992 800 261112
rect 289451 256504 290251 256624
rect 0 253920 800 254040
rect 289451 249976 290251 250096
rect 0 246984 800 247104
rect 289451 243448 290251 243568
rect 0 240048 800 240168
rect 289451 237056 290251 237176
rect 0 233112 800 233232
rect 289451 230528 290251 230648
rect 0 226176 800 226296
rect 289451 224000 290251 224120
rect 0 219104 800 219224
rect 289451 217472 290251 217592
rect 0 212168 800 212288
rect 289451 210944 290251 211064
rect 0 205232 800 205352
rect 289451 204552 290251 204672
rect 0 198296 800 198416
rect 289451 198024 290251 198144
rect 0 191360 800 191480
rect 289451 191496 290251 191616
rect 289451 184968 290251 185088
rect 0 184288 800 184408
rect 289451 178576 290251 178696
rect 0 177352 800 177472
rect 289451 172048 290251 172168
rect 0 170416 800 170536
rect 289451 165520 290251 165640
rect 0 163480 800 163600
rect 289451 158992 290251 159112
rect 0 156544 800 156664
rect 289451 152464 290251 152584
rect 0 149608 800 149728
rect 289451 146072 290251 146192
rect 0 142536 800 142656
rect 289451 139544 290251 139664
rect 0 135600 800 135720
rect 289451 133016 290251 133136
rect 0 128664 800 128784
rect 289451 126488 290251 126608
rect 0 121728 800 121848
rect 289451 120096 290251 120216
rect 0 114792 800 114912
rect 289451 113568 290251 113688
rect 0 107720 800 107840
rect 289451 107040 290251 107160
rect 0 100784 800 100904
rect 289451 100512 290251 100632
rect 0 93848 800 93968
rect 289451 93984 290251 94104
rect 289451 87592 290251 87712
rect 0 86912 800 87032
rect 289451 81064 290251 81184
rect 0 79976 800 80096
rect 289451 74536 290251 74656
rect 0 72904 800 73024
rect 289451 68008 290251 68128
rect 0 65968 800 66088
rect 289451 61616 290251 61736
rect 0 59032 800 59152
rect 289451 55088 290251 55208
rect 0 52096 800 52216
rect 289451 48560 290251 48680
rect 0 45160 800 45280
rect 289451 42032 290251 42152
rect 0 38088 800 38208
rect 289451 35504 290251 35624
rect 0 31152 800 31272
rect 289451 29112 290251 29232
rect 0 24216 800 24336
rect 289451 22584 290251 22704
rect 0 17280 800 17400
rect 289451 16056 290251 16176
rect 0 10344 800 10464
rect 289451 9528 290251 9648
rect 0 3408 800 3528
rect 289451 3136 290251 3256
<< obsm3 >>
rect 289 289208 289451 289985
rect 289 288936 289371 289208
rect 880 288928 289371 288936
rect 880 288656 289451 288928
rect 289 282680 289451 288656
rect 289 282400 289371 282680
rect 289 282000 289451 282400
rect 880 281720 289451 282000
rect 289 276152 289451 281720
rect 289 275872 289371 276152
rect 289 275064 289451 275872
rect 880 274784 289451 275064
rect 289 269624 289451 274784
rect 289 269344 289371 269624
rect 289 268128 289451 269344
rect 880 267848 289451 268128
rect 289 263232 289451 267848
rect 289 262952 289371 263232
rect 289 261192 289451 262952
rect 880 260912 289451 261192
rect 289 256704 289451 260912
rect 289 256424 289371 256704
rect 289 254120 289451 256424
rect 880 253840 289451 254120
rect 289 250176 289451 253840
rect 289 249896 289371 250176
rect 289 247184 289451 249896
rect 880 246904 289451 247184
rect 289 243648 289451 246904
rect 289 243368 289371 243648
rect 289 240248 289451 243368
rect 880 239968 289451 240248
rect 289 237256 289451 239968
rect 289 236976 289371 237256
rect 289 233312 289451 236976
rect 880 233032 289451 233312
rect 289 230728 289451 233032
rect 289 230448 289371 230728
rect 289 226376 289451 230448
rect 880 226096 289451 226376
rect 289 224200 289451 226096
rect 289 223920 289371 224200
rect 289 219304 289451 223920
rect 880 219024 289451 219304
rect 289 217672 289451 219024
rect 289 217392 289371 217672
rect 289 212368 289451 217392
rect 880 212088 289451 212368
rect 289 211144 289451 212088
rect 289 210864 289371 211144
rect 289 205432 289451 210864
rect 880 205152 289451 205432
rect 289 204752 289451 205152
rect 289 204472 289371 204752
rect 289 198496 289451 204472
rect 880 198224 289451 198496
rect 880 198216 289371 198224
rect 289 197944 289371 198216
rect 289 191696 289451 197944
rect 289 191560 289371 191696
rect 880 191416 289371 191560
rect 880 191280 289451 191416
rect 289 185168 289451 191280
rect 289 184888 289371 185168
rect 289 184488 289451 184888
rect 880 184208 289451 184488
rect 289 178776 289451 184208
rect 289 178496 289371 178776
rect 289 177552 289451 178496
rect 880 177272 289451 177552
rect 289 172248 289451 177272
rect 289 171968 289371 172248
rect 289 170616 289451 171968
rect 880 170336 289451 170616
rect 289 165720 289451 170336
rect 289 165440 289371 165720
rect 289 163680 289451 165440
rect 880 163400 289451 163680
rect 289 159192 289451 163400
rect 289 158912 289371 159192
rect 289 156744 289451 158912
rect 880 156464 289451 156744
rect 289 152664 289451 156464
rect 289 152384 289371 152664
rect 289 149808 289451 152384
rect 880 149528 289451 149808
rect 289 146272 289451 149528
rect 289 145992 289371 146272
rect 289 142736 289451 145992
rect 880 142456 289451 142736
rect 289 139744 289451 142456
rect 289 139464 289371 139744
rect 289 135800 289451 139464
rect 880 135520 289451 135800
rect 289 133216 289451 135520
rect 289 132936 289371 133216
rect 289 128864 289451 132936
rect 880 128584 289451 128864
rect 289 126688 289451 128584
rect 289 126408 289371 126688
rect 289 121928 289451 126408
rect 880 121648 289451 121928
rect 289 120296 289451 121648
rect 289 120016 289371 120296
rect 289 114992 289451 120016
rect 880 114712 289451 114992
rect 289 113768 289451 114712
rect 289 113488 289371 113768
rect 289 107920 289451 113488
rect 880 107640 289451 107920
rect 289 107240 289451 107640
rect 289 106960 289371 107240
rect 289 100984 289451 106960
rect 880 100712 289451 100984
rect 880 100704 289371 100712
rect 289 100432 289371 100704
rect 289 94184 289451 100432
rect 289 94048 289371 94184
rect 880 93904 289371 94048
rect 880 93768 289451 93904
rect 289 87792 289451 93768
rect 289 87512 289371 87792
rect 289 87112 289451 87512
rect 880 86832 289451 87112
rect 289 81264 289451 86832
rect 289 80984 289371 81264
rect 289 80176 289451 80984
rect 880 79896 289451 80176
rect 289 74736 289451 79896
rect 289 74456 289371 74736
rect 289 73104 289451 74456
rect 880 72824 289451 73104
rect 289 68208 289451 72824
rect 289 67928 289371 68208
rect 289 66168 289451 67928
rect 880 65888 289451 66168
rect 289 61816 289451 65888
rect 289 61536 289371 61816
rect 289 59232 289451 61536
rect 880 58952 289451 59232
rect 289 55288 289451 58952
rect 289 55008 289371 55288
rect 289 52296 289451 55008
rect 880 52016 289451 52296
rect 289 48760 289451 52016
rect 289 48480 289371 48760
rect 289 45360 289451 48480
rect 880 45080 289451 45360
rect 289 42232 289451 45080
rect 289 41952 289371 42232
rect 289 38288 289451 41952
rect 880 38008 289451 38288
rect 289 35704 289451 38008
rect 289 35424 289371 35704
rect 289 31352 289451 35424
rect 880 31072 289451 31352
rect 289 29312 289451 31072
rect 289 29032 289371 29312
rect 289 24416 289451 29032
rect 880 24136 289451 24416
rect 289 22784 289451 24136
rect 289 22504 289371 22784
rect 289 17480 289451 22504
rect 880 17200 289451 17480
rect 289 16256 289451 17200
rect 289 15976 289371 16256
rect 289 10544 289451 15976
rect 880 10264 289451 10544
rect 289 9728 289451 10264
rect 289 9448 289371 9728
rect 289 3608 289451 9448
rect 880 3336 289451 3608
rect 880 3328 289371 3336
rect 289 3056 289371 3328
rect 289 851 289451 3056
<< metal4 >>
rect 4208 2128 4528 290000
rect 4868 2176 5188 289952
rect 5528 2176 5848 289952
rect 6188 2176 6508 289952
rect 19568 2128 19888 290000
rect 20228 2176 20548 289952
rect 20888 2176 21208 289952
rect 21548 2176 21868 289952
rect 34928 2128 35248 290000
rect 35588 2176 35908 289952
rect 36248 2176 36568 289952
rect 36908 2176 37228 289952
rect 50288 2128 50608 290000
rect 50948 2176 51268 289952
rect 51608 2176 51928 289952
rect 52268 2176 52588 289952
rect 65648 2128 65968 290000
rect 66308 2176 66628 289952
rect 66968 2176 67288 289952
rect 67628 2176 67948 289952
rect 81008 2128 81328 290000
rect 81668 2176 81988 289952
rect 82328 2176 82648 289952
rect 82988 2176 83308 289952
rect 96368 2128 96688 290000
rect 97028 2176 97348 289952
rect 97688 2176 98008 289952
rect 98348 2176 98668 289952
rect 111728 2128 112048 290000
rect 112388 2176 112708 289952
rect 113048 2176 113368 289952
rect 113708 2176 114028 289952
rect 127088 2128 127408 290000
rect 127748 2176 128068 289952
rect 128408 2176 128728 289952
rect 129068 2176 129388 289952
rect 142448 2128 142768 290000
rect 143108 2176 143428 289952
rect 143768 2176 144088 289952
rect 144428 2176 144748 289952
rect 157808 2128 158128 290000
rect 158468 2176 158788 289952
rect 159128 2176 159448 289952
rect 159788 2176 160108 289952
rect 173168 2128 173488 290000
rect 173828 2176 174148 289952
rect 174488 2176 174808 289952
rect 175148 2176 175468 289952
rect 188528 2128 188848 290000
rect 189188 2176 189508 289952
rect 189848 2176 190168 289952
rect 190508 2176 190828 289952
rect 203888 2128 204208 290000
rect 204548 2176 204868 289952
rect 205208 2176 205528 289952
rect 205868 2176 206188 289952
rect 219248 2128 219568 290000
rect 219908 2176 220228 289952
rect 220568 2176 220888 289952
rect 221228 2176 221548 289952
rect 234608 2128 234928 290000
rect 235268 2176 235588 289952
rect 235928 2176 236248 289952
rect 236588 2176 236908 289952
rect 249968 2128 250288 290000
rect 250628 2176 250948 289952
rect 251288 2176 251608 289952
rect 251948 2176 252268 289952
rect 265328 2128 265648 290000
rect 265988 2176 266308 289952
rect 266648 2176 266968 289952
rect 267308 2176 267628 289952
rect 280688 2128 281008 290000
rect 281348 2176 281668 289952
rect 282008 2176 282328 289952
rect 282668 2176 282988 289952
<< obsm4 >>
rect 3739 2619 4128 255101
rect 4608 2619 4788 255101
rect 5268 2619 5448 255101
rect 5928 2619 6108 255101
rect 6588 2619 19488 255101
rect 19968 2619 20148 255101
rect 20628 2619 20808 255101
rect 21288 2619 21468 255101
rect 21948 2619 34848 255101
rect 35328 2619 35508 255101
rect 35988 2619 36168 255101
rect 36648 2619 36828 255101
rect 37308 2619 50208 255101
rect 50688 2619 50868 255101
rect 51348 2619 51528 255101
rect 52008 2619 52188 255101
rect 52668 2619 65568 255101
rect 66048 2619 66228 255101
rect 66708 2619 66888 255101
rect 67368 2619 67548 255101
rect 68028 2619 80928 255101
rect 81408 2619 81588 255101
rect 82068 2619 82248 255101
rect 82728 2619 82908 255101
rect 83388 2619 96288 255101
rect 96768 2619 96948 255101
rect 97428 2619 97608 255101
rect 98088 2619 98268 255101
rect 98748 2619 111648 255101
rect 112128 2619 112308 255101
rect 112788 2619 112968 255101
rect 113448 2619 113628 255101
rect 114108 2619 127008 255101
rect 127488 2619 127668 255101
rect 128148 2619 128328 255101
rect 128808 2619 128988 255101
rect 129468 2619 142368 255101
rect 142848 2619 143028 255101
rect 143508 2619 143688 255101
rect 144168 2619 144348 255101
rect 144828 2619 157728 255101
rect 158208 2619 158388 255101
rect 158868 2619 159048 255101
rect 159528 2619 159708 255101
rect 160188 2619 173088 255101
rect 173568 2619 173748 255101
rect 174228 2619 174408 255101
rect 174888 2619 175068 255101
rect 175548 2619 188448 255101
rect 188928 2619 189108 255101
rect 189588 2619 189768 255101
rect 190248 2619 190428 255101
rect 190908 2619 203808 255101
rect 204288 2619 204468 255101
rect 204948 2619 205128 255101
rect 205608 2619 205788 255101
rect 206268 2619 219168 255101
rect 219648 2619 219828 255101
rect 220308 2619 220488 255101
rect 220968 2619 221148 255101
rect 221628 2619 234528 255101
rect 235008 2619 235188 255101
rect 235668 2619 235848 255101
rect 236328 2619 236508 255101
rect 236988 2619 249888 255101
rect 250368 2619 250548 255101
rect 251028 2619 251208 255101
rect 251688 2619 251837 255101
<< labels >>
rlabel metal3 s 289451 3136 290251 3256 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 289451 198024 290251 198144 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 289451 217472 290251 217592 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 289451 237056 290251 237176 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 289451 256504 290251 256624 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 289451 275952 290251 276072 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 284850 291595 284906 292395 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 252558 291595 252614 292395 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 220358 291595 220414 292395 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 188066 291595 188122 292395 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 155774 291595 155830 292395 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 289451 22584 290251 22704 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 123574 291595 123630 292395 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 91282 291595 91338 292395 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 59082 291595 59138 292395 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 26790 291595 26846 292395 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 274864 800 274984 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 253920 800 254040 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 233112 800 233232 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 212168 800 212288 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 191360 800 191480 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 170416 800 170536 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 289451 42032 290251 42152 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 149608 800 149728 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 128664 800 128784 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 107720 800 107840 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 86912 800 87032 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 65968 800 66088 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 45160 800 45280 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 289451 61616 290251 61736 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 289451 81064 290251 81184 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 289451 100512 290251 100632 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 289451 120096 290251 120216 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 289451 139544 290251 139664 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 289451 158992 290251 159112 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 289451 178576 290251 178696 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 289451 16056 290251 16176 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 289451 210944 290251 211064 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 289451 230528 290251 230648 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 289451 249976 290251 250096 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 289451 269424 290251 269544 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 289451 289008 290251 289128 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 263322 291595 263378 292395 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 231030 291595 231086 292395 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 198830 291595 198886 292395 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 166538 291595 166594 292395 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 134338 291595 134394 292395 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 289451 35504 290251 35624 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 102046 291595 102102 292395 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 69846 291595 69902 292395 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 37554 291595 37610 292395 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 5354 291595 5410 292395 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 288736 800 288856 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 267928 800 268048 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 246984 800 247104 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 226176 800 226296 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 205232 800 205352 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 184288 800 184408 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 289451 55088 290251 55208 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 163480 800 163600 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 142536 800 142656 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 121728 800 121848 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 100784 800 100904 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 79976 800 80096 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 59032 800 59152 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 17280 800 17400 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 289451 74536 290251 74656 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 289451 93984 290251 94104 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 289451 113568 290251 113688 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 289451 133016 290251 133136 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 289451 152464 290251 152584 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 289451 172048 290251 172168 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 289451 191496 290251 191616 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 289451 9528 290251 9648 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 289451 204552 290251 204672 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 289451 224000 290251 224120 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 289451 243448 290251 243568 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 289451 263032 290251 263152 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 289451 282480 290251 282600 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 274086 291595 274142 292395 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 241794 291595 241850 292395 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 209594 291595 209650 292395 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 177302 291595 177358 292395 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 145102 291595 145158 292395 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 289451 29112 290251 29232 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 112810 291595 112866 292395 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 80518 291595 80574 292395 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 48318 291595 48374 292395 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 16026 291595 16082 292395 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 281800 800 281920 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 260992 800 261112 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 240048 800 240168 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 219104 800 219224 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 198296 800 198416 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 177352 800 177472 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 289451 48560 290251 48680 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 156544 800 156664 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 135600 800 135720 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 114792 800 114912 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 93848 800 93968 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 72904 800 73024 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 52096 800 52216 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 31152 800 31272 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 289451 68008 290251 68128 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 289451 87592 290251 87712 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 289451 107040 290251 107160 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 289451 126488 290251 126608 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 289451 146072 290251 146192 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 289451 165520 290251 165640 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 289451 184968 290251 185088 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 240782 0 240838 800 6 la_data_in[100]
port 116 nsew signal input
rlabel metal2 s 242530 0 242586 800 6 la_data_in[101]
port 117 nsew signal input
rlabel metal2 s 244278 0 244334 800 6 la_data_in[102]
port 118 nsew signal input
rlabel metal2 s 246118 0 246174 800 6 la_data_in[103]
port 119 nsew signal input
rlabel metal2 s 247866 0 247922 800 6 la_data_in[104]
port 120 nsew signal input
rlabel metal2 s 249614 0 249670 800 6 la_data_in[105]
port 121 nsew signal input
rlabel metal2 s 251454 0 251510 800 6 la_data_in[106]
port 122 nsew signal input
rlabel metal2 s 253202 0 253258 800 6 la_data_in[107]
port 123 nsew signal input
rlabel metal2 s 254950 0 255006 800 6 la_data_in[108]
port 124 nsew signal input
rlabel metal2 s 256698 0 256754 800 6 la_data_in[109]
port 125 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_data_in[10]
port 126 nsew signal input
rlabel metal2 s 258538 0 258594 800 6 la_data_in[110]
port 127 nsew signal input
rlabel metal2 s 260286 0 260342 800 6 la_data_in[111]
port 128 nsew signal input
rlabel metal2 s 262034 0 262090 800 6 la_data_in[112]
port 129 nsew signal input
rlabel metal2 s 263874 0 263930 800 6 la_data_in[113]
port 130 nsew signal input
rlabel metal2 s 265622 0 265678 800 6 la_data_in[114]
port 131 nsew signal input
rlabel metal2 s 267370 0 267426 800 6 la_data_in[115]
port 132 nsew signal input
rlabel metal2 s 269210 0 269266 800 6 la_data_in[116]
port 133 nsew signal input
rlabel metal2 s 270958 0 271014 800 6 la_data_in[117]
port 134 nsew signal input
rlabel metal2 s 272706 0 272762 800 6 la_data_in[118]
port 135 nsew signal input
rlabel metal2 s 274546 0 274602 800 6 la_data_in[119]
port 136 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_data_in[11]
port 137 nsew signal input
rlabel metal2 s 276294 0 276350 800 6 la_data_in[120]
port 138 nsew signal input
rlabel metal2 s 278042 0 278098 800 6 la_data_in[121]
port 139 nsew signal input
rlabel metal2 s 279882 0 279938 800 6 la_data_in[122]
port 140 nsew signal input
rlabel metal2 s 281630 0 281686 800 6 la_data_in[123]
port 141 nsew signal input
rlabel metal2 s 283378 0 283434 800 6 la_data_in[124]
port 142 nsew signal input
rlabel metal2 s 285218 0 285274 800 6 la_data_in[125]
port 143 nsew signal input
rlabel metal2 s 286966 0 287022 800 6 la_data_in[126]
port 144 nsew signal input
rlabel metal2 s 288714 0 288770 800 6 la_data_in[127]
port 145 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_data_in[12]
port 146 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_data_in[13]
port 147 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_data_in[14]
port 148 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_data_in[15]
port 149 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 la_data_in[16]
port 150 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_data_in[17]
port 151 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 la_data_in[18]
port 152 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_data_in[19]
port 153 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 la_data_in[1]
port 154 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_data_in[20]
port 155 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_data_in[21]
port 156 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 la_data_in[22]
port 157 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 la_data_in[23]
port 158 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 la_data_in[24]
port 159 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 la_data_in[25]
port 160 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 la_data_in[26]
port 161 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 la_data_in[27]
port 162 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 la_data_in[28]
port 163 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 la_data_in[29]
port 164 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_data_in[2]
port 165 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_data_in[30]
port 166 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_data_in[31]
port 167 nsew signal input
rlabel metal2 s 119894 0 119950 800 6 la_data_in[32]
port 168 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 la_data_in[33]
port 169 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 la_data_in[34]
port 170 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 la_data_in[35]
port 171 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_data_in[36]
port 172 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 la_data_in[37]
port 173 nsew signal input
rlabel metal2 s 130566 0 130622 800 6 la_data_in[38]
port 174 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 la_data_in[39]
port 175 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_data_in[3]
port 176 nsew signal input
rlabel metal2 s 134154 0 134210 800 6 la_data_in[40]
port 177 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_data_in[41]
port 178 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 la_data_in[42]
port 179 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 la_data_in[43]
port 180 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 la_data_in[44]
port 181 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 la_data_in[45]
port 182 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 la_data_in[46]
port 183 nsew signal input
rlabel metal2 s 146574 0 146630 800 6 la_data_in[47]
port 184 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 la_data_in[48]
port 185 nsew signal input
rlabel metal2 s 150162 0 150218 800 6 la_data_in[49]
port 186 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_data_in[4]
port 187 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 la_data_in[50]
port 188 nsew signal input
rlabel metal2 s 153658 0 153714 800 6 la_data_in[51]
port 189 nsew signal input
rlabel metal2 s 155406 0 155462 800 6 la_data_in[52]
port 190 nsew signal input
rlabel metal2 s 157246 0 157302 800 6 la_data_in[53]
port 191 nsew signal input
rlabel metal2 s 158994 0 159050 800 6 la_data_in[54]
port 192 nsew signal input
rlabel metal2 s 160742 0 160798 800 6 la_data_in[55]
port 193 nsew signal input
rlabel metal2 s 162582 0 162638 800 6 la_data_in[56]
port 194 nsew signal input
rlabel metal2 s 164330 0 164386 800 6 la_data_in[57]
port 195 nsew signal input
rlabel metal2 s 166078 0 166134 800 6 la_data_in[58]
port 196 nsew signal input
rlabel metal2 s 167918 0 167974 800 6 la_data_in[59]
port 197 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_data_in[5]
port 198 nsew signal input
rlabel metal2 s 169666 0 169722 800 6 la_data_in[60]
port 199 nsew signal input
rlabel metal2 s 171414 0 171470 800 6 la_data_in[61]
port 200 nsew signal input
rlabel metal2 s 173254 0 173310 800 6 la_data_in[62]
port 201 nsew signal input
rlabel metal2 s 175002 0 175058 800 6 la_data_in[63]
port 202 nsew signal input
rlabel metal2 s 176750 0 176806 800 6 la_data_in[64]
port 203 nsew signal input
rlabel metal2 s 178590 0 178646 800 6 la_data_in[65]
port 204 nsew signal input
rlabel metal2 s 180338 0 180394 800 6 la_data_in[66]
port 205 nsew signal input
rlabel metal2 s 182086 0 182142 800 6 la_data_in[67]
port 206 nsew signal input
rlabel metal2 s 183926 0 183982 800 6 la_data_in[68]
port 207 nsew signal input
rlabel metal2 s 185674 0 185730 800 6 la_data_in[69]
port 208 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_data_in[6]
port 209 nsew signal input
rlabel metal2 s 187422 0 187478 800 6 la_data_in[70]
port 210 nsew signal input
rlabel metal2 s 189170 0 189226 800 6 la_data_in[71]
port 211 nsew signal input
rlabel metal2 s 191010 0 191066 800 6 la_data_in[72]
port 212 nsew signal input
rlabel metal2 s 192758 0 192814 800 6 la_data_in[73]
port 213 nsew signal input
rlabel metal2 s 194506 0 194562 800 6 la_data_in[74]
port 214 nsew signal input
rlabel metal2 s 196346 0 196402 800 6 la_data_in[75]
port 215 nsew signal input
rlabel metal2 s 198094 0 198150 800 6 la_data_in[76]
port 216 nsew signal input
rlabel metal2 s 199842 0 199898 800 6 la_data_in[77]
port 217 nsew signal input
rlabel metal2 s 201682 0 201738 800 6 la_data_in[78]
port 218 nsew signal input
rlabel metal2 s 203430 0 203486 800 6 la_data_in[79]
port 219 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_data_in[7]
port 220 nsew signal input
rlabel metal2 s 205178 0 205234 800 6 la_data_in[80]
port 221 nsew signal input
rlabel metal2 s 207018 0 207074 800 6 la_data_in[81]
port 222 nsew signal input
rlabel metal2 s 208766 0 208822 800 6 la_data_in[82]
port 223 nsew signal input
rlabel metal2 s 210514 0 210570 800 6 la_data_in[83]
port 224 nsew signal input
rlabel metal2 s 212354 0 212410 800 6 la_data_in[84]
port 225 nsew signal input
rlabel metal2 s 214102 0 214158 800 6 la_data_in[85]
port 226 nsew signal input
rlabel metal2 s 215850 0 215906 800 6 la_data_in[86]
port 227 nsew signal input
rlabel metal2 s 217690 0 217746 800 6 la_data_in[87]
port 228 nsew signal input
rlabel metal2 s 219438 0 219494 800 6 la_data_in[88]
port 229 nsew signal input
rlabel metal2 s 221186 0 221242 800 6 la_data_in[89]
port 230 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la_data_in[8]
port 231 nsew signal input
rlabel metal2 s 222934 0 222990 800 6 la_data_in[90]
port 232 nsew signal input
rlabel metal2 s 224774 0 224830 800 6 la_data_in[91]
port 233 nsew signal input
rlabel metal2 s 226522 0 226578 800 6 la_data_in[92]
port 234 nsew signal input
rlabel metal2 s 228270 0 228326 800 6 la_data_in[93]
port 235 nsew signal input
rlabel metal2 s 230110 0 230166 800 6 la_data_in[94]
port 236 nsew signal input
rlabel metal2 s 231858 0 231914 800 6 la_data_in[95]
port 237 nsew signal input
rlabel metal2 s 233606 0 233662 800 6 la_data_in[96]
port 238 nsew signal input
rlabel metal2 s 235446 0 235502 800 6 la_data_in[97]
port 239 nsew signal input
rlabel metal2 s 237194 0 237250 800 6 la_data_in[98]
port 240 nsew signal input
rlabel metal2 s 238942 0 238998 800 6 la_data_in[99]
port 241 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_data_in[9]
port 242 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_data_out[0]
port 243 nsew signal output
rlabel metal2 s 241334 0 241390 800 6 la_data_out[100]
port 244 nsew signal output
rlabel metal2 s 243082 0 243138 800 6 la_data_out[101]
port 245 nsew signal output
rlabel metal2 s 244922 0 244978 800 6 la_data_out[102]
port 246 nsew signal output
rlabel metal2 s 246670 0 246726 800 6 la_data_out[103]
port 247 nsew signal output
rlabel metal2 s 248418 0 248474 800 6 la_data_out[104]
port 248 nsew signal output
rlabel metal2 s 250258 0 250314 800 6 la_data_out[105]
port 249 nsew signal output
rlabel metal2 s 252006 0 252062 800 6 la_data_out[106]
port 250 nsew signal output
rlabel metal2 s 253754 0 253810 800 6 la_data_out[107]
port 251 nsew signal output
rlabel metal2 s 255594 0 255650 800 6 la_data_out[108]
port 252 nsew signal output
rlabel metal2 s 257342 0 257398 800 6 la_data_out[109]
port 253 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 la_data_out[10]
port 254 nsew signal output
rlabel metal2 s 259090 0 259146 800 6 la_data_out[110]
port 255 nsew signal output
rlabel metal2 s 260930 0 260986 800 6 la_data_out[111]
port 256 nsew signal output
rlabel metal2 s 262678 0 262734 800 6 la_data_out[112]
port 257 nsew signal output
rlabel metal2 s 264426 0 264482 800 6 la_data_out[113]
port 258 nsew signal output
rlabel metal2 s 266266 0 266322 800 6 la_data_out[114]
port 259 nsew signal output
rlabel metal2 s 268014 0 268070 800 6 la_data_out[115]
port 260 nsew signal output
rlabel metal2 s 269762 0 269818 800 6 la_data_out[116]
port 261 nsew signal output
rlabel metal2 s 271510 0 271566 800 6 la_data_out[117]
port 262 nsew signal output
rlabel metal2 s 273350 0 273406 800 6 la_data_out[118]
port 263 nsew signal output
rlabel metal2 s 275098 0 275154 800 6 la_data_out[119]
port 264 nsew signal output
rlabel metal2 s 83186 0 83242 800 6 la_data_out[11]
port 265 nsew signal output
rlabel metal2 s 276846 0 276902 800 6 la_data_out[120]
port 266 nsew signal output
rlabel metal2 s 278686 0 278742 800 6 la_data_out[121]
port 267 nsew signal output
rlabel metal2 s 280434 0 280490 800 6 la_data_out[122]
port 268 nsew signal output
rlabel metal2 s 282182 0 282238 800 6 la_data_out[123]
port 269 nsew signal output
rlabel metal2 s 284022 0 284078 800 6 la_data_out[124]
port 270 nsew signal output
rlabel metal2 s 285770 0 285826 800 6 la_data_out[125]
port 271 nsew signal output
rlabel metal2 s 287518 0 287574 800 6 la_data_out[126]
port 272 nsew signal output
rlabel metal2 s 289358 0 289414 800 6 la_data_out[127]
port 273 nsew signal output
rlabel metal2 s 84934 0 84990 800 6 la_data_out[12]
port 274 nsew signal output
rlabel metal2 s 86774 0 86830 800 6 la_data_out[13]
port 275 nsew signal output
rlabel metal2 s 88522 0 88578 800 6 la_data_out[14]
port 276 nsew signal output
rlabel metal2 s 90270 0 90326 800 6 la_data_out[15]
port 277 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 la_data_out[16]
port 278 nsew signal output
rlabel metal2 s 93858 0 93914 800 6 la_data_out[17]
port 279 nsew signal output
rlabel metal2 s 95606 0 95662 800 6 la_data_out[18]
port 280 nsew signal output
rlabel metal2 s 97354 0 97410 800 6 la_data_out[19]
port 281 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 la_data_out[1]
port 282 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 la_data_out[20]
port 283 nsew signal output
rlabel metal2 s 100942 0 100998 800 6 la_data_out[21]
port 284 nsew signal output
rlabel metal2 s 102690 0 102746 800 6 la_data_out[22]
port 285 nsew signal output
rlabel metal2 s 104530 0 104586 800 6 la_data_out[23]
port 286 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 la_data_out[24]
port 287 nsew signal output
rlabel metal2 s 108026 0 108082 800 6 la_data_out[25]
port 288 nsew signal output
rlabel metal2 s 109866 0 109922 800 6 la_data_out[26]
port 289 nsew signal output
rlabel metal2 s 111614 0 111670 800 6 la_data_out[27]
port 290 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 la_data_out[28]
port 291 nsew signal output
rlabel metal2 s 115202 0 115258 800 6 la_data_out[29]
port 292 nsew signal output
rlabel metal2 s 67178 0 67234 800 6 la_data_out[2]
port 293 nsew signal output
rlabel metal2 s 116950 0 117006 800 6 la_data_out[30]
port 294 nsew signal output
rlabel metal2 s 118698 0 118754 800 6 la_data_out[31]
port 295 nsew signal output
rlabel metal2 s 120538 0 120594 800 6 la_data_out[32]
port 296 nsew signal output
rlabel metal2 s 122286 0 122342 800 6 la_data_out[33]
port 297 nsew signal output
rlabel metal2 s 124034 0 124090 800 6 la_data_out[34]
port 298 nsew signal output
rlabel metal2 s 125874 0 125930 800 6 la_data_out[35]
port 299 nsew signal output
rlabel metal2 s 127622 0 127678 800 6 la_data_out[36]
port 300 nsew signal output
rlabel metal2 s 129370 0 129426 800 6 la_data_out[37]
port 301 nsew signal output
rlabel metal2 s 131118 0 131174 800 6 la_data_out[38]
port 302 nsew signal output
rlabel metal2 s 132958 0 133014 800 6 la_data_out[39]
port 303 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 la_data_out[3]
port 304 nsew signal output
rlabel metal2 s 134706 0 134762 800 6 la_data_out[40]
port 305 nsew signal output
rlabel metal2 s 136454 0 136510 800 6 la_data_out[41]
port 306 nsew signal output
rlabel metal2 s 138294 0 138350 800 6 la_data_out[42]
port 307 nsew signal output
rlabel metal2 s 140042 0 140098 800 6 la_data_out[43]
port 308 nsew signal output
rlabel metal2 s 141790 0 141846 800 6 la_data_out[44]
port 309 nsew signal output
rlabel metal2 s 143630 0 143686 800 6 la_data_out[45]
port 310 nsew signal output
rlabel metal2 s 145378 0 145434 800 6 la_data_out[46]
port 311 nsew signal output
rlabel metal2 s 147126 0 147182 800 6 la_data_out[47]
port 312 nsew signal output
rlabel metal2 s 148966 0 149022 800 6 la_data_out[48]
port 313 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 la_data_out[49]
port 314 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 la_data_out[4]
port 315 nsew signal output
rlabel metal2 s 152462 0 152518 800 6 la_data_out[50]
port 316 nsew signal output
rlabel metal2 s 154302 0 154358 800 6 la_data_out[51]
port 317 nsew signal output
rlabel metal2 s 156050 0 156106 800 6 la_data_out[52]
port 318 nsew signal output
rlabel metal2 s 157798 0 157854 800 6 la_data_out[53]
port 319 nsew signal output
rlabel metal2 s 159638 0 159694 800 6 la_data_out[54]
port 320 nsew signal output
rlabel metal2 s 161386 0 161442 800 6 la_data_out[55]
port 321 nsew signal output
rlabel metal2 s 163134 0 163190 800 6 la_data_out[56]
port 322 nsew signal output
rlabel metal2 s 164882 0 164938 800 6 la_data_out[57]
port 323 nsew signal output
rlabel metal2 s 166722 0 166778 800 6 la_data_out[58]
port 324 nsew signal output
rlabel metal2 s 168470 0 168526 800 6 la_data_out[59]
port 325 nsew signal output
rlabel metal2 s 72514 0 72570 800 6 la_data_out[5]
port 326 nsew signal output
rlabel metal2 s 170218 0 170274 800 6 la_data_out[60]
port 327 nsew signal output
rlabel metal2 s 172058 0 172114 800 6 la_data_out[61]
port 328 nsew signal output
rlabel metal2 s 173806 0 173862 800 6 la_data_out[62]
port 329 nsew signal output
rlabel metal2 s 175554 0 175610 800 6 la_data_out[63]
port 330 nsew signal output
rlabel metal2 s 177394 0 177450 800 6 la_data_out[64]
port 331 nsew signal output
rlabel metal2 s 179142 0 179198 800 6 la_data_out[65]
port 332 nsew signal output
rlabel metal2 s 180890 0 180946 800 6 la_data_out[66]
port 333 nsew signal output
rlabel metal2 s 182730 0 182786 800 6 la_data_out[67]
port 334 nsew signal output
rlabel metal2 s 184478 0 184534 800 6 la_data_out[68]
port 335 nsew signal output
rlabel metal2 s 186226 0 186282 800 6 la_data_out[69]
port 336 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 la_data_out[6]
port 337 nsew signal output
rlabel metal2 s 188066 0 188122 800 6 la_data_out[70]
port 338 nsew signal output
rlabel metal2 s 189814 0 189870 800 6 la_data_out[71]
port 339 nsew signal output
rlabel metal2 s 191562 0 191618 800 6 la_data_out[72]
port 340 nsew signal output
rlabel metal2 s 193402 0 193458 800 6 la_data_out[73]
port 341 nsew signal output
rlabel metal2 s 195150 0 195206 800 6 la_data_out[74]
port 342 nsew signal output
rlabel metal2 s 196898 0 196954 800 6 la_data_out[75]
port 343 nsew signal output
rlabel metal2 s 198646 0 198702 800 6 la_data_out[76]
port 344 nsew signal output
rlabel metal2 s 200486 0 200542 800 6 la_data_out[77]
port 345 nsew signal output
rlabel metal2 s 202234 0 202290 800 6 la_data_out[78]
port 346 nsew signal output
rlabel metal2 s 203982 0 204038 800 6 la_data_out[79]
port 347 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 la_data_out[7]
port 348 nsew signal output
rlabel metal2 s 205822 0 205878 800 6 la_data_out[80]
port 349 nsew signal output
rlabel metal2 s 207570 0 207626 800 6 la_data_out[81]
port 350 nsew signal output
rlabel metal2 s 209318 0 209374 800 6 la_data_out[82]
port 351 nsew signal output
rlabel metal2 s 211158 0 211214 800 6 la_data_out[83]
port 352 nsew signal output
rlabel metal2 s 212906 0 212962 800 6 la_data_out[84]
port 353 nsew signal output
rlabel metal2 s 214654 0 214710 800 6 la_data_out[85]
port 354 nsew signal output
rlabel metal2 s 216494 0 216550 800 6 la_data_out[86]
port 355 nsew signal output
rlabel metal2 s 218242 0 218298 800 6 la_data_out[87]
port 356 nsew signal output
rlabel metal2 s 219990 0 220046 800 6 la_data_out[88]
port 357 nsew signal output
rlabel metal2 s 221830 0 221886 800 6 la_data_out[89]
port 358 nsew signal output
rlabel metal2 s 77850 0 77906 800 6 la_data_out[8]
port 359 nsew signal output
rlabel metal2 s 223578 0 223634 800 6 la_data_out[90]
port 360 nsew signal output
rlabel metal2 s 225326 0 225382 800 6 la_data_out[91]
port 361 nsew signal output
rlabel metal2 s 227166 0 227222 800 6 la_data_out[92]
port 362 nsew signal output
rlabel metal2 s 228914 0 228970 800 6 la_data_out[93]
port 363 nsew signal output
rlabel metal2 s 230662 0 230718 800 6 la_data_out[94]
port 364 nsew signal output
rlabel metal2 s 232502 0 232558 800 6 la_data_out[95]
port 365 nsew signal output
rlabel metal2 s 234250 0 234306 800 6 la_data_out[96]
port 366 nsew signal output
rlabel metal2 s 235998 0 236054 800 6 la_data_out[97]
port 367 nsew signal output
rlabel metal2 s 237746 0 237802 800 6 la_data_out[98]
port 368 nsew signal output
rlabel metal2 s 239586 0 239642 800 6 la_data_out[99]
port 369 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 la_data_out[9]
port 370 nsew signal output
rlabel metal2 s 64234 0 64290 800 6 la_oen[0]
port 371 nsew signal input
rlabel metal2 s 241978 0 242034 800 6 la_oen[100]
port 372 nsew signal input
rlabel metal2 s 243726 0 243782 800 6 la_oen[101]
port 373 nsew signal input
rlabel metal2 s 245474 0 245530 800 6 la_oen[102]
port 374 nsew signal input
rlabel metal2 s 247222 0 247278 800 6 la_oen[103]
port 375 nsew signal input
rlabel metal2 s 249062 0 249118 800 6 la_oen[104]
port 376 nsew signal input
rlabel metal2 s 250810 0 250866 800 6 la_oen[105]
port 377 nsew signal input
rlabel metal2 s 252558 0 252614 800 6 la_oen[106]
port 378 nsew signal input
rlabel metal2 s 254398 0 254454 800 6 la_oen[107]
port 379 nsew signal input
rlabel metal2 s 256146 0 256202 800 6 la_oen[108]
port 380 nsew signal input
rlabel metal2 s 257894 0 257950 800 6 la_oen[109]
port 381 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_oen[10]
port 382 nsew signal input
rlabel metal2 s 259734 0 259790 800 6 la_oen[110]
port 383 nsew signal input
rlabel metal2 s 261482 0 261538 800 6 la_oen[111]
port 384 nsew signal input
rlabel metal2 s 263230 0 263286 800 6 la_oen[112]
port 385 nsew signal input
rlabel metal2 s 265070 0 265126 800 6 la_oen[113]
port 386 nsew signal input
rlabel metal2 s 266818 0 266874 800 6 la_oen[114]
port 387 nsew signal input
rlabel metal2 s 268566 0 268622 800 6 la_oen[115]
port 388 nsew signal input
rlabel metal2 s 270406 0 270462 800 6 la_oen[116]
port 389 nsew signal input
rlabel metal2 s 272154 0 272210 800 6 la_oen[117]
port 390 nsew signal input
rlabel metal2 s 273902 0 273958 800 6 la_oen[118]
port 391 nsew signal input
rlabel metal2 s 275742 0 275798 800 6 la_oen[119]
port 392 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_oen[11]
port 393 nsew signal input
rlabel metal2 s 277490 0 277546 800 6 la_oen[120]
port 394 nsew signal input
rlabel metal2 s 279238 0 279294 800 6 la_oen[121]
port 395 nsew signal input
rlabel metal2 s 280986 0 281042 800 6 la_oen[122]
port 396 nsew signal input
rlabel metal2 s 282826 0 282882 800 6 la_oen[123]
port 397 nsew signal input
rlabel metal2 s 284574 0 284630 800 6 la_oen[124]
port 398 nsew signal input
rlabel metal2 s 286322 0 286378 800 6 la_oen[125]
port 399 nsew signal input
rlabel metal2 s 288162 0 288218 800 6 la_oen[126]
port 400 nsew signal input
rlabel metal2 s 289910 0 289966 800 6 la_oen[127]
port 401 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 la_oen[12]
port 402 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_oen[13]
port 403 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_oen[14]
port 404 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_oen[15]
port 405 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_oen[16]
port 406 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 la_oen[17]
port 407 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_oen[18]
port 408 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_oen[19]
port 409 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_oen[1]
port 410 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_oen[20]
port 411 nsew signal input
rlabel metal2 s 101586 0 101642 800 6 la_oen[21]
port 412 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 la_oen[22]
port 413 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 la_oen[23]
port 414 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 la_oen[24]
port 415 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 la_oen[25]
port 416 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 la_oen[26]
port 417 nsew signal input
rlabel metal2 s 112166 0 112222 800 6 la_oen[27]
port 418 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_oen[28]
port 419 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 la_oen[29]
port 420 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_oen[2]
port 421 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 la_oen[30]
port 422 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 la_oen[31]
port 423 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 la_oen[32]
port 424 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 la_oen[33]
port 425 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 la_oen[34]
port 426 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 la_oen[35]
port 427 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 la_oen[36]
port 428 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 la_oen[37]
port 429 nsew signal input
rlabel metal2 s 131762 0 131818 800 6 la_oen[38]
port 430 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 la_oen[39]
port 431 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_oen[3]
port 432 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 la_oen[40]
port 433 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 la_oen[41]
port 434 nsew signal input
rlabel metal2 s 138846 0 138902 800 6 la_oen[42]
port 435 nsew signal input
rlabel metal2 s 140594 0 140650 800 6 la_oen[43]
port 436 nsew signal input
rlabel metal2 s 142434 0 142490 800 6 la_oen[44]
port 437 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_oen[45]
port 438 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 la_oen[46]
port 439 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_oen[47]
port 440 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 la_oen[48]
port 441 nsew signal input
rlabel metal2 s 151266 0 151322 800 6 la_oen[49]
port 442 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_oen[4]
port 443 nsew signal input
rlabel metal2 s 153106 0 153162 800 6 la_oen[50]
port 444 nsew signal input
rlabel metal2 s 154854 0 154910 800 6 la_oen[51]
port 445 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_oen[52]
port 446 nsew signal input
rlabel metal2 s 158442 0 158498 800 6 la_oen[53]
port 447 nsew signal input
rlabel metal2 s 160190 0 160246 800 6 la_oen[54]
port 448 nsew signal input
rlabel metal2 s 161938 0 161994 800 6 la_oen[55]
port 449 nsew signal input
rlabel metal2 s 163778 0 163834 800 6 la_oen[56]
port 450 nsew signal input
rlabel metal2 s 165526 0 165582 800 6 la_oen[57]
port 451 nsew signal input
rlabel metal2 s 167274 0 167330 800 6 la_oen[58]
port 452 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 la_oen[59]
port 453 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_oen[5]
port 454 nsew signal input
rlabel metal2 s 170862 0 170918 800 6 la_oen[60]
port 455 nsew signal input
rlabel metal2 s 172610 0 172666 800 6 la_oen[61]
port 456 nsew signal input
rlabel metal2 s 174450 0 174506 800 6 la_oen[62]
port 457 nsew signal input
rlabel metal2 s 176198 0 176254 800 6 la_oen[63]
port 458 nsew signal input
rlabel metal2 s 177946 0 178002 800 6 la_oen[64]
port 459 nsew signal input
rlabel metal2 s 179694 0 179750 800 6 la_oen[65]
port 460 nsew signal input
rlabel metal2 s 181534 0 181590 800 6 la_oen[66]
port 461 nsew signal input
rlabel metal2 s 183282 0 183338 800 6 la_oen[67]
port 462 nsew signal input
rlabel metal2 s 185030 0 185086 800 6 la_oen[68]
port 463 nsew signal input
rlabel metal2 s 186870 0 186926 800 6 la_oen[69]
port 464 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 la_oen[6]
port 465 nsew signal input
rlabel metal2 s 188618 0 188674 800 6 la_oen[70]
port 466 nsew signal input
rlabel metal2 s 190366 0 190422 800 6 la_oen[71]
port 467 nsew signal input
rlabel metal2 s 192206 0 192262 800 6 la_oen[72]
port 468 nsew signal input
rlabel metal2 s 193954 0 194010 800 6 la_oen[73]
port 469 nsew signal input
rlabel metal2 s 195702 0 195758 800 6 la_oen[74]
port 470 nsew signal input
rlabel metal2 s 197542 0 197598 800 6 la_oen[75]
port 471 nsew signal input
rlabel metal2 s 199290 0 199346 800 6 la_oen[76]
port 472 nsew signal input
rlabel metal2 s 201038 0 201094 800 6 la_oen[77]
port 473 nsew signal input
rlabel metal2 s 202878 0 202934 800 6 la_oen[78]
port 474 nsew signal input
rlabel metal2 s 204626 0 204682 800 6 la_oen[79]
port 475 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_oen[7]
port 476 nsew signal input
rlabel metal2 s 206374 0 206430 800 6 la_oen[80]
port 477 nsew signal input
rlabel metal2 s 208214 0 208270 800 6 la_oen[81]
port 478 nsew signal input
rlabel metal2 s 209962 0 210018 800 6 la_oen[82]
port 479 nsew signal input
rlabel metal2 s 211710 0 211766 800 6 la_oen[83]
port 480 nsew signal input
rlabel metal2 s 213458 0 213514 800 6 la_oen[84]
port 481 nsew signal input
rlabel metal2 s 215298 0 215354 800 6 la_oen[85]
port 482 nsew signal input
rlabel metal2 s 217046 0 217102 800 6 la_oen[86]
port 483 nsew signal input
rlabel metal2 s 218794 0 218850 800 6 la_oen[87]
port 484 nsew signal input
rlabel metal2 s 220634 0 220690 800 6 la_oen[88]
port 485 nsew signal input
rlabel metal2 s 222382 0 222438 800 6 la_oen[89]
port 486 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_oen[8]
port 487 nsew signal input
rlabel metal2 s 224130 0 224186 800 6 la_oen[90]
port 488 nsew signal input
rlabel metal2 s 225970 0 226026 800 6 la_oen[91]
port 489 nsew signal input
rlabel metal2 s 227718 0 227774 800 6 la_oen[92]
port 490 nsew signal input
rlabel metal2 s 229466 0 229522 800 6 la_oen[93]
port 491 nsew signal input
rlabel metal2 s 231306 0 231362 800 6 la_oen[94]
port 492 nsew signal input
rlabel metal2 s 233054 0 233110 800 6 la_oen[95]
port 493 nsew signal input
rlabel metal2 s 234802 0 234858 800 6 la_oen[96]
port 494 nsew signal input
rlabel metal2 s 236642 0 236698 800 6 la_oen[97]
port 495 nsew signal input
rlabel metal2 s 238390 0 238446 800 6 la_oen[98]
port 496 nsew signal input
rlabel metal2 s 240138 0 240194 800 6 la_oen[99]
port 497 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 la_oen[9]
port 498 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 499 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_rst_i
port 500 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_ack_o
port 501 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 wbs_adr_i[0]
port 502 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_adr_i[10]
port 503 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_adr_i[11]
port 504 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_adr_i[12]
port 505 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_adr_i[13]
port 506 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_adr_i[14]
port 507 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wbs_adr_i[15]
port 508 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 wbs_adr_i[16]
port 509 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_adr_i[17]
port 510 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wbs_adr_i[18]
port 511 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 wbs_adr_i[19]
port 512 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_adr_i[1]
port 513 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 wbs_adr_i[20]
port 514 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 wbs_adr_i[21]
port 515 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 wbs_adr_i[22]
port 516 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 wbs_adr_i[23]
port 517 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 wbs_adr_i[24]
port 518 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 wbs_adr_i[25]
port 519 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 wbs_adr_i[26]
port 520 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 wbs_adr_i[27]
port 521 nsew signal input
rlabel metal2 s 55954 0 56010 800 6 wbs_adr_i[28]
port 522 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 wbs_adr_i[29]
port 523 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_adr_i[2]
port 524 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 wbs_adr_i[30]
port 525 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 wbs_adr_i[31]
port 526 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_adr_i[3]
port 527 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_adr_i[4]
port 528 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_adr_i[5]
port 529 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_adr_i[6]
port 530 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_adr_i[7]
port 531 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[8]
port 532 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_adr_i[9]
port 533 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_cyc_i
port 534 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_i[0]
port 535 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_dat_i[10]
port 536 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_dat_i[11]
port 537 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_i[12]
port 538 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 wbs_dat_i[13]
port 539 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 wbs_dat_i[14]
port 540 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wbs_dat_i[15]
port 541 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 wbs_dat_i[16]
port 542 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 wbs_dat_i[17]
port 543 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 wbs_dat_i[18]
port 544 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wbs_dat_i[19]
port 545 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_i[1]
port 546 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 wbs_dat_i[20]
port 547 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 wbs_dat_i[21]
port 548 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 wbs_dat_i[22]
port 549 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 wbs_dat_i[23]
port 550 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 wbs_dat_i[24]
port 551 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 wbs_dat_i[25]
port 552 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 wbs_dat_i[26]
port 553 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 wbs_dat_i[27]
port 554 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 wbs_dat_i[28]
port 555 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 wbs_dat_i[29]
port 556 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_dat_i[2]
port 557 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 wbs_dat_i[30]
port 558 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 wbs_dat_i[31]
port 559 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_i[3]
port 560 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_i[4]
port 561 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_i[5]
port 562 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_i[6]
port 563 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_i[7]
port 564 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_i[8]
port 565 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_dat_i[9]
port 566 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_dat_o[0]
port 567 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_o[10]
port 568 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_o[11]
port 569 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_o[12]
port 570 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_o[13]
port 571 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_o[14]
port 572 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 wbs_dat_o[15]
port 573 nsew signal output
rlabel metal2 s 35806 0 35862 800 6 wbs_dat_o[16]
port 574 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 wbs_dat_o[17]
port 575 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 wbs_dat_o[18]
port 576 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 wbs_dat_o[19]
port 577 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[1]
port 578 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 wbs_dat_o[20]
port 579 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 wbs_dat_o[21]
port 580 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 wbs_dat_o[22]
port 581 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 wbs_dat_o[23]
port 582 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 wbs_dat_o[24]
port 583 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 wbs_dat_o[25]
port 584 nsew signal output
rlabel metal2 s 53562 0 53618 800 6 wbs_dat_o[26]
port 585 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 wbs_dat_o[27]
port 586 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 wbs_dat_o[28]
port 587 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 wbs_dat_o[29]
port 588 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[2]
port 589 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 wbs_dat_o[30]
port 590 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 wbs_dat_o[31]
port 591 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_o[3]
port 592 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_o[4]
port 593 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_o[5]
port 594 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_o[6]
port 595 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_o[7]
port 596 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_o[8]
port 597 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_o[9]
port 598 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 wbs_sel_i[0]
port 599 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_sel_i[1]
port 600 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_sel_i[2]
port 601 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_sel_i[3]
port 602 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_stb_i
port 603 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_we_i
port 604 nsew signal input
rlabel metal4 s 280688 2128 281008 290000 6 vccd1
port 605 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 290000 6 vccd1
port 606 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 290000 6 vccd1
port 607 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 290000 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 290000 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 290000 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 290000 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 290000 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 290000 6 vccd1
port 613 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 290000 6 vccd1
port 614 nsew power bidirectional
rlabel metal4 s 265328 2128 265648 290000 6 vssd1
port 615 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 290000 6 vssd1
port 616 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 290000 6 vssd1
port 617 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 290000 6 vssd1
port 618 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 290000 6 vssd1
port 619 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 290000 6 vssd1
port 620 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 290000 6 vssd1
port 621 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 290000 6 vssd1
port 622 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 290000 6 vssd1
port 623 nsew ground bidirectional
rlabel metal4 s 281348 2176 281668 289952 6 vccd2
port 624 nsew power bidirectional
rlabel metal4 s 250628 2176 250948 289952 6 vccd2
port 625 nsew power bidirectional
rlabel metal4 s 219908 2176 220228 289952 6 vccd2
port 626 nsew power bidirectional
rlabel metal4 s 189188 2176 189508 289952 6 vccd2
port 627 nsew power bidirectional
rlabel metal4 s 158468 2176 158788 289952 6 vccd2
port 628 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 289952 6 vccd2
port 629 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 289952 6 vccd2
port 630 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 289952 6 vccd2
port 631 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 289952 6 vccd2
port 632 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 289952 6 vccd2
port 633 nsew power bidirectional
rlabel metal4 s 265988 2176 266308 289952 6 vssd2
port 634 nsew ground bidirectional
rlabel metal4 s 235268 2176 235588 289952 6 vssd2
port 635 nsew ground bidirectional
rlabel metal4 s 204548 2176 204868 289952 6 vssd2
port 636 nsew ground bidirectional
rlabel metal4 s 173828 2176 174148 289952 6 vssd2
port 637 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 289952 6 vssd2
port 638 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 289952 6 vssd2
port 639 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 289952 6 vssd2
port 640 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 289952 6 vssd2
port 641 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 289952 6 vssd2
port 642 nsew ground bidirectional
rlabel metal4 s 282008 2176 282328 289952 6 vdda1
port 643 nsew power bidirectional
rlabel metal4 s 251288 2176 251608 289952 6 vdda1
port 644 nsew power bidirectional
rlabel metal4 s 220568 2176 220888 289952 6 vdda1
port 645 nsew power bidirectional
rlabel metal4 s 189848 2176 190168 289952 6 vdda1
port 646 nsew power bidirectional
rlabel metal4 s 159128 2176 159448 289952 6 vdda1
port 647 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 289952 6 vdda1
port 648 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 289952 6 vdda1
port 649 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 289952 6 vdda1
port 650 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 289952 6 vdda1
port 651 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 289952 6 vdda1
port 652 nsew power bidirectional
rlabel metal4 s 266648 2176 266968 289952 6 vssa1
port 653 nsew ground bidirectional
rlabel metal4 s 235928 2176 236248 289952 6 vssa1
port 654 nsew ground bidirectional
rlabel metal4 s 205208 2176 205528 289952 6 vssa1
port 655 nsew ground bidirectional
rlabel metal4 s 174488 2176 174808 289952 6 vssa1
port 656 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 289952 6 vssa1
port 657 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 289952 6 vssa1
port 658 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 289952 6 vssa1
port 659 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 289952 6 vssa1
port 660 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 289952 6 vssa1
port 661 nsew ground bidirectional
rlabel metal4 s 282668 2176 282988 289952 6 vdda2
port 662 nsew power bidirectional
rlabel metal4 s 251948 2176 252268 289952 6 vdda2
port 663 nsew power bidirectional
rlabel metal4 s 221228 2176 221548 289952 6 vdda2
port 664 nsew power bidirectional
rlabel metal4 s 190508 2176 190828 289952 6 vdda2
port 665 nsew power bidirectional
rlabel metal4 s 159788 2176 160108 289952 6 vdda2
port 666 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 289952 6 vdda2
port 667 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 289952 6 vdda2
port 668 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 289952 6 vdda2
port 669 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 289952 6 vdda2
port 670 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 289952 6 vdda2
port 671 nsew power bidirectional
rlabel metal4 s 267308 2176 267628 289952 6 vssa2
port 672 nsew ground bidirectional
rlabel metal4 s 236588 2176 236908 289952 6 vssa2
port 673 nsew ground bidirectional
rlabel metal4 s 205868 2176 206188 289952 6 vssa2
port 674 nsew ground bidirectional
rlabel metal4 s 175148 2176 175468 289952 6 vssa2
port 675 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 289952 6 vssa2
port 676 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 289952 6 vssa2
port 677 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 289952 6 vssa2
port 678 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 289952 6 vssa2
port 679 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 289952 6 vssa2
port 680 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 290251 292395
string LEFview TRUE
<< end >>

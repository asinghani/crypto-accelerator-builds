* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for accelerator_top abstract view
.subckt accelerator_top io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oen[0] la_oen[100] la_oen[101]
+ la_oen[102] la_oen[103] la_oen[104] la_oen[105] la_oen[106] la_oen[107] la_oen[108]
+ la_oen[109] la_oen[10] la_oen[110] la_oen[111] la_oen[112] la_oen[113] la_oen[114]
+ la_oen[115] la_oen[116] la_oen[117] la_oen[118] la_oen[119] la_oen[11] la_oen[120]
+ la_oen[121] la_oen[122] la_oen[123] la_oen[124] la_oen[125] la_oen[126] la_oen[127]
+ la_oen[12] la_oen[13] la_oen[14] la_oen[15] la_oen[16] la_oen[17] la_oen[18] la_oen[19]
+ la_oen[1] la_oen[20] la_oen[21] la_oen[22] la_oen[23] la_oen[24] la_oen[25] la_oen[26]
+ la_oen[27] la_oen[28] la_oen[29] la_oen[2] la_oen[30] la_oen[31] la_oen[32] la_oen[33]
+ la_oen[34] la_oen[35] la_oen[36] la_oen[37] la_oen[38] la_oen[39] la_oen[3] la_oen[40]
+ la_oen[41] la_oen[42] la_oen[43] la_oen[44] la_oen[45] la_oen[46] la_oen[47] la_oen[48]
+ la_oen[49] la_oen[4] la_oen[50] la_oen[51] la_oen[52] la_oen[53] la_oen[54] la_oen[55]
+ la_oen[56] la_oen[57] la_oen[58] la_oen[59] la_oen[5] la_oen[60] la_oen[61] la_oen[62]
+ la_oen[63] la_oen[64] la_oen[65] la_oen[66] la_oen[67] la_oen[68] la_oen[69] la_oen[6]
+ la_oen[70] la_oen[71] la_oen[72] la_oen[73] la_oen[74] la_oen[75] la_oen[76] la_oen[77]
+ la_oen[78] la_oen[79] la_oen[7] la_oen[80] la_oen[81] la_oen[82] la_oen[83] la_oen[84]
+ la_oen[85] la_oen[86] la_oen[87] la_oen[88] la_oen[89] la_oen[8] la_oen[90] la_oen[91]
+ la_oen[92] la_oen[93] la_oen[94] la_oen[95] la_oen[96] la_oen[97] la_oen[98] la_oen[99]
+ la_oen[9] wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i VPWR VGND
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[29]
+ analog_io[2] analog_io[30] analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7]
+ analog_io[8] analog_io[9] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oen[0] la_oen[100] la_oen[101]
+ la_oen[102] la_oen[103] la_oen[104] la_oen[105] la_oen[106] la_oen[107] la_oen[108]
+ la_oen[109] la_oen[10] la_oen[110] la_oen[111] la_oen[112] la_oen[113] la_oen[114]
+ la_oen[115] la_oen[116] la_oen[117] la_oen[118] la_oen[119] la_oen[11] la_oen[120]
+ la_oen[121] la_oen[122] la_oen[123] la_oen[124] la_oen[125] la_oen[126] la_oen[127]
+ la_oen[12] la_oen[13] la_oen[14] la_oen[15] la_oen[16] la_oen[17] la_oen[18] la_oen[19]
+ la_oen[1] la_oen[20] la_oen[21] la_oen[22] la_oen[23] la_oen[24] la_oen[25] la_oen[26]
+ la_oen[27] la_oen[28] la_oen[29] la_oen[2] la_oen[30] la_oen[31] la_oen[32] la_oen[33]
+ la_oen[34] la_oen[35] la_oen[36] la_oen[37] la_oen[38] la_oen[39] la_oen[3] la_oen[40]
+ la_oen[41] la_oen[42] la_oen[43] la_oen[44] la_oen[45] la_oen[46] la_oen[47] la_oen[48]
+ la_oen[49] la_oen[4] la_oen[50] la_oen[51] la_oen[52] la_oen[53] la_oen[54] la_oen[55]
+ la_oen[56] la_oen[57] la_oen[58] la_oen[59] la_oen[5] la_oen[60] la_oen[61] la_oen[62]
+ la_oen[63] la_oen[64] la_oen[65] la_oen[66] la_oen[67] la_oen[68] la_oen[69] la_oen[6]
+ la_oen[70] la_oen[71] la_oen[72] la_oen[73] la_oen[74] la_oen[75] la_oen[76] la_oen[77]
+ la_oen[78] la_oen[79] la_oen[7] la_oen[80] la_oen[81] la_oen[82] la_oen[83] la_oen[84]
+ la_oen[85] la_oen[86] la_oen[87] la_oen[88] la_oen[89] la_oen[8] la_oen[90] la_oen[91]
+ la_oen[92] la_oen[93] la_oen[94] la_oen[95] la_oen[96] la_oen[97] la_oen[98] la_oen[99]
+ la_oen[9] user_clock2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
+ vccd1 vssd1 vccd2 vssd2 vdda1 vssa1 vdda2 vssa2
XANTENNA_mprj_la_oen[125] la_oen[125] ANTENNA_mprj_la_oen[125]/VGND VSUBS ANTENNA_mprj_la_oen[125]/VPB
+ ANTENNA_mprj_la_oen[125]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[100] la_data_in[100] ANTENNA_mprj_la_data_in[100]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[100]/VPB ANTENNA_mprj_la_data_in[100]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[13] la_data_in[13] ANTENNA_mprj_la_data_in[13]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[13]/VPB ANTENNA_mprj_la_data_in[13]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[10] wbs_adr_i[10] ANTENNA_mprj_wbs_adr_i[10]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[10]/VPB
+ ANTENNA_mprj_wbs_adr_i[10]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[23] wbs_dat_i[23] ANTENNA_mprj_wbs_dat_i[23]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[23]/VPB
+ ANTENNA_mprj_wbs_dat_i[23]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[5] la_oen[5] ANTENNA_mprj_la_oen[5]/VGND VSUBS ANTENNA_mprj_la_oen[5]/VPB
+ ANTENNA_mprj_la_oen[5]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[108] la_oen[108] ANTENNA_mprj_la_oen[108]/VGND VSUBS ANTENNA_mprj_la_oen[108]/VPB
+ ANTENNA_mprj_la_oen[108]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[82] la_oen[82] ANTENNA_mprj_la_oen[82]/VGND VSUBS ANTENNA_mprj_la_oen[82]/VPB
+ ANTENNA_mprj_la_oen[82]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[65] la_oen[65] ANTENNA_mprj_la_oen[65]/VGND VSUBS ANTENNA_mprj_la_oen[65]/VPB
+ ANTENNA_mprj_la_oen[65]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[2] wbs_dat_i[2] ANTENNA_mprj_wbs_dat_i[2]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[2]/VPB
+ ANTENNA_mprj_wbs_dat_i[2]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[48] la_oen[48] ANTENNA_mprj_la_oen[48]/VGND VSUBS ANTENNA_mprj_la_oen[48]/VPB
+ ANTENNA_mprj_la_oen[48]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[1] wbs_adr_i[1] ANTENNA_mprj_wbs_adr_i[1]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[1]/VPB
+ ANTENNA_mprj_wbs_adr_i[1]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_sel_i[2] wbs_sel_i[2] ANTENNA_mprj_wbs_sel_i[2]/VGND VSUBS ANTENNA_mprj_wbs_sel_i[2]/VPB
+ ANTENNA_mprj_wbs_sel_i[2]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[89] la_data_in[89] ANTENNA_mprj_la_data_in[89]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[89]/VPB ANTENNA_mprj_la_data_in[89]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[12] la_data_in[12] ANTENNA_mprj_la_data_in[12]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[12]/VPB ANTENNA_mprj_la_data_in[12]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[124] la_oen[124] ANTENNA_mprj_la_oen[124]/VGND VSUBS ANTENNA_mprj_la_oen[124]/VPB
+ ANTENNA_mprj_la_oen[124]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[81] la_oen[81] ANTENNA_mprj_la_oen[81]/VGND VSUBS ANTENNA_mprj_la_oen[81]/VPB
+ ANTENNA_mprj_la_oen[81]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[22] wbs_dat_i[22] ANTENNA_mprj_wbs_dat_i[22]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[22]/VPB
+ ANTENNA_mprj_wbs_dat_i[22]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[4] la_oen[4] ANTENNA_mprj_la_oen[4]/VGND VSUBS ANTENNA_mprj_la_oen[4]/VPB
+ ANTENNA_mprj_la_oen[4]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[107] la_oen[107] ANTENNA_mprj_la_oen[107]/VGND VSUBS ANTENNA_mprj_la_oen[107]/VPB
+ ANTENNA_mprj_la_oen[107]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[64] la_oen[64] ANTENNA_mprj_la_oen[64]/VGND VSUBS ANTENNA_mprj_la_oen[64]/VPB
+ ANTENNA_mprj_la_oen[64]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[0] wbs_adr_i[0] ANTENNA_mprj_wbs_adr_i[0]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[0]/VPB
+ ANTENNA_mprj_wbs_adr_i[0]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[1] wbs_dat_i[1] ANTENNA_mprj_wbs_dat_i[1]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[1]/VPB
+ ANTENNA_mprj_wbs_dat_i[1]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_sel_i[1] wbs_sel_i[1] ANTENNA_mprj_wbs_sel_i[1]/VGND VSUBS ANTENNA_mprj_wbs_sel_i[1]/VPB
+ ANTENNA_mprj_wbs_sel_i[1]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[47] la_oen[47] ANTENNA_mprj_la_oen[47]/VGND VSUBS ANTENNA_mprj_la_oen[47]/VPB
+ ANTENNA_mprj_la_oen[47]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[123] la_oen[123] ANTENNA_mprj_la_oen[123]/VGND VSUBS ANTENNA_mprj_la_oen[123]/VPB
+ ANTENNA_mprj_la_oen[123]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[88] la_data_in[88] ANTENNA_mprj_la_data_in[88]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[88]/VPB ANTENNA_mprj_la_data_in[88]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[21] wbs_dat_i[21] ANTENNA_mprj_wbs_dat_i[21]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[21]/VPB
+ ANTENNA_mprj_wbs_dat_i[21]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[3] la_oen[3] ANTENNA_mprj_la_oen[3]/VGND VSUBS ANTENNA_mprj_la_oen[3]/VPB
+ ANTENNA_mprj_la_oen[3]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[11] la_data_in[11] ANTENNA_mprj_la_data_in[11]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[11]/VPB ANTENNA_mprj_la_data_in[11]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[106] la_oen[106] ANTENNA_mprj_la_oen[106]/VGND VSUBS ANTENNA_mprj_la_oen[106]/VPB
+ ANTENNA_mprj_la_oen[106]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[80] la_oen[80] ANTENNA_mprj_la_oen[80]/VGND VSUBS ANTENNA_mprj_la_oen[80]/VPB
+ ANTENNA_mprj_la_oen[80]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[0] wbs_dat_i[0] ANTENNA_mprj_wbs_dat_i[0]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[0]/VPB
+ ANTENNA_mprj_wbs_dat_i[0]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[63] la_oen[63] ANTENNA_mprj_la_oen[63]/VGND VSUBS ANTENNA_mprj_la_oen[63]/VPB
+ ANTENNA_mprj_la_oen[63]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[46] la_oen[46] ANTENNA_mprj_la_oen[46]/VGND VSUBS ANTENNA_mprj_la_oen[46]/VPB
+ ANTENNA_mprj_la_oen[46]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_sel_i[0] wbs_sel_i[0] ANTENNA_mprj_wbs_sel_i[0]/VGND VSUBS ANTENNA_mprj_wbs_sel_i[0]/VPB
+ ANTENNA_mprj_wbs_sel_i[0]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[87] la_data_in[87] ANTENNA_mprj_la_data_in[87]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[87]/VPB ANTENNA_mprj_la_data_in[87]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[29] la_oen[29] ANTENNA_mprj_la_oen[29]/VGND VSUBS ANTENNA_mprj_la_oen[29]/VPB
+ ANTENNA_mprj_la_oen[29]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[122] la_oen[122] ANTENNA_mprj_la_oen[122]/VGND VSUBS ANTENNA_mprj_la_oen[122]/VPB
+ ANTENNA_mprj_la_oen[122]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[20] wbs_dat_i[20] ANTENNA_mprj_wbs_dat_i[20]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[20]/VPB
+ ANTENNA_mprj_wbs_dat_i[20]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[2] la_oen[2] ANTENNA_mprj_la_oen[2]/VGND VSUBS ANTENNA_mprj_la_oen[2]/VPB
+ ANTENNA_mprj_la_oen[2]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[10] la_data_in[10] ANTENNA_mprj_la_data_in[10]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[10]/VPB ANTENNA_mprj_la_data_in[10]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[105] la_oen[105] ANTENNA_mprj_la_oen[105]/VGND VSUBS ANTENNA_mprj_la_oen[105]/VPB
+ ANTENNA_mprj_la_oen[105]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[62] la_oen[62] ANTENNA_mprj_la_oen[62]/VGND VSUBS ANTENNA_mprj_la_oen[62]/VPB
+ ANTENNA_mprj_la_oen[62]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[45] la_oen[45] ANTENNA_mprj_la_oen[45]/VGND VSUBS ANTENNA_mprj_la_oen[45]/VPB
+ ANTENNA_mprj_la_oen[45]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[28] la_oen[28] ANTENNA_mprj_la_oen[28]/VGND VSUBS ANTENNA_mprj_la_oen[28]/VPB
+ ANTENNA_mprj_la_oen[28]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[29] io_in[29] ANTENNA_mprj_io_in[29]/VGND VSUBS ANTENNA_mprj_io_in[29]/VPB
+ ANTENNA_mprj_io_in[29]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[86] la_data_in[86] ANTENNA_mprj_la_data_in[86]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[86]/VPB ANTENNA_mprj_la_data_in[86]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[69] la_data_in[69] ANTENNA_mprj_la_data_in[69]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[69]/VPB ANTENNA_mprj_la_data_in[69]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[1] la_oen[1] ANTENNA_mprj_la_oen[1]/VGND VSUBS ANTENNA_mprj_la_oen[1]/VPB
+ ANTENNA_mprj_la_oen[1]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[121] la_oen[121] ANTENNA_mprj_la_oen[121]/VGND VSUBS ANTENNA_mprj_la_oen[121]/VPB
+ ANTENNA_mprj_la_oen[121]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[104] la_oen[104] ANTENNA_mprj_la_oen[104]/VGND VSUBS ANTENNA_mprj_la_oen[104]/VPB
+ ANTENNA_mprj_la_oen[104]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[61] la_oen[61] ANTENNA_mprj_la_oen[61]/VGND VSUBS ANTENNA_mprj_la_oen[61]/VPB
+ ANTENNA_mprj_la_oen[61]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[44] la_oen[44] ANTENNA_mprj_la_oen[44]/VGND VSUBS ANTENNA_mprj_la_oen[44]/VPB
+ ANTENNA_mprj_la_oen[44]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[28] io_in[28] ANTENNA_mprj_io_in[28]/VGND VSUBS ANTENNA_mprj_io_in[28]/VPB
+ ANTENNA_mprj_io_in[28]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[85] la_data_in[85] ANTENNA_mprj_la_data_in[85]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[85]/VPB ANTENNA_mprj_la_data_in[85]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[27] la_oen[27] ANTENNA_mprj_la_oen[27]/VGND VSUBS ANTENNA_mprj_la_oen[27]/VPB
+ ANTENNA_mprj_la_oen[27]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[120] la_oen[120] ANTENNA_mprj_la_oen[120]/VGND VSUBS ANTENNA_mprj_la_oen[120]/VPB
+ ANTENNA_mprj_la_oen[120]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[68] la_data_in[68] ANTENNA_mprj_la_data_in[68]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[68]/VPB ANTENNA_mprj_la_data_in[68]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[0] la_oen[0] ANTENNA_mprj_la_oen[0]/VGND VSUBS ANTENNA_mprj_la_oen[0]/VPB
+ ANTENNA_mprj_la_oen[0]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[103] la_oen[103] ANTENNA_mprj_la_oen[103]/VGND VSUBS ANTENNA_mprj_la_oen[103]/VPB
+ ANTENNA_mprj_la_oen[103]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[60] la_oen[60] ANTENNA_mprj_la_oen[60]/VGND VSUBS ANTENNA_mprj_la_oen[60]/VPB
+ ANTENNA_mprj_la_oen[60]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[43] la_oen[43] ANTENNA_mprj_la_oen[43]/VGND VSUBS ANTENNA_mprj_la_oen[43]/VPB
+ ANTENNA_mprj_la_oen[43]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[26] la_oen[26] ANTENNA_mprj_la_oen[26]/VGND VSUBS ANTENNA_mprj_la_oen[26]/VPB
+ ANTENNA_mprj_la_oen[26]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[27] io_in[27] ANTENNA_mprj_io_in[27]/VGND VSUBS ANTENNA_mprj_io_in[27]/VPB
+ ANTENNA_mprj_io_in[27]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[84] la_data_in[84] ANTENNA_mprj_la_data_in[84]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[84]/VPB ANTENNA_mprj_la_data_in[84]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[67] la_data_in[67] ANTENNA_mprj_la_data_in[67]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[67]/VPB ANTENNA_mprj_la_data_in[67]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[102] la_oen[102] ANTENNA_mprj_la_oen[102]/VGND VSUBS ANTENNA_mprj_la_oen[102]/VPB
+ ANTENNA_mprj_la_oen[102]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[42] la_oen[42] ANTENNA_mprj_la_oen[42]/VGND VSUBS ANTENNA_mprj_la_oen[42]/VPB
+ ANTENNA_mprj_la_oen[42]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[26] io_in[26] ANTENNA_mprj_io_in[26]/VGND VSUBS ANTENNA_mprj_io_in[26]/VPB
+ ANTENNA_mprj_io_in[26]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[83] la_data_in[83] ANTENNA_mprj_la_data_in[83]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[83]/VPB ANTENNA_mprj_la_data_in[83]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[25] la_oen[25] ANTENNA_mprj_la_oen[25]/VGND VSUBS ANTENNA_mprj_la_oen[25]/VPB
+ ANTENNA_mprj_la_oen[25]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wb_rst_i wb_rst_i ANTENNA_mprj_wb_clk_i/VGND VSUBS ANTENNA_mprj_wb_rst_i/VPB
+ ANTENNA_mprj_wb_rst_i/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[66] la_data_in[66] ANTENNA_mprj_la_data_in[66]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[66]/VPB ANTENNA_mprj_la_data_in[66]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[119] la_data_in[119] ANTENNA_mprj_la_data_in[119]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[119]/VPB ANTENNA_mprj_la_data_in[119]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[101] la_oen[101] ANTENNA_mprj_la_oen[101]/VGND VSUBS ANTENNA_mprj_la_oen[101]/VPB
+ ANTENNA_mprj_la_oen[101]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[49] la_data_in[49] ANTENNA_mprj_la_data_in[49]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[49]/VPB ANTENNA_mprj_la_data_in[49]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[41] la_oen[41] ANTENNA_mprj_la_oen[41]/VGND VSUBS ANTENNA_mprj_la_oen[41]/VPB
+ ANTENNA_mprj_la_oen[41]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[29] wbs_adr_i[29] ANTENNA_mprj_wbs_adr_i[29]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[29]/VPB
+ ANTENNA_mprj_wbs_adr_i[29]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[25] io_in[25] ANTENNA_mprj_io_in[25]/VGND VSUBS ANTENNA_mprj_io_in[25]/VPB
+ ANTENNA_mprj_io_in[25]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[82] la_data_in[82] ANTENNA_mprj_la_data_in[82]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[82]/VPB ANTENNA_mprj_la_data_in[82]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[24] la_oen[24] ANTENNA_mprj_la_oen[24]/VGND VSUBS ANTENNA_mprj_la_oen[24]/VPB
+ ANTENNA_mprj_la_oen[24]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[100] la_oen[100] ANTENNA_mprj_la_oen[100]/VGND VSUBS ANTENNA_mprj_la_oen[100]/VPB
+ ANTENNA_mprj_la_oen[100]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[65] la_data_in[65] ANTENNA_mprj_la_data_in[65]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[65]/VPB ANTENNA_mprj_la_data_in[65]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[48] la_data_in[48] ANTENNA_mprj_la_data_in[48]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[48]/VPB ANTENNA_mprj_la_data_in[48]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[118] la_data_in[118] ANTENNA_mprj_la_data_in[118]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[118]/VPB ANTENNA_mprj_la_data_in[118]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[40] la_oen[40] ANTENNA_mprj_la_oen[40]/VGND VSUBS ANTENNA_mprj_la_oen[40]/VPB
+ ANTENNA_mprj_la_oen[40]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[28] wbs_adr_i[28] ANTENNA_mprj_wbs_adr_i[28]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[28]/VPB
+ ANTENNA_mprj_wbs_adr_i[28]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[24] io_in[24] ANTENNA_mprj_io_in[24]/VGND VSUBS ANTENNA_mprj_io_in[24]/VPB
+ ANTENNA_mprj_io_in[24]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[81] la_data_in[81] ANTENNA_mprj_la_data_in[81]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[81]/VPB ANTENNA_mprj_la_data_in[81]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[23] la_oen[23] ANTENNA_mprj_la_oen[23]/VGND VSUBS ANTENNA_mprj_la_oen[23]/VPB
+ ANTENNA_mprj_la_oen[23]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[64] la_data_in[64] ANTENNA_mprj_la_data_in[64]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[64]/VPB ANTENNA_mprj_la_data_in[64]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[117] la_data_in[117] ANTENNA_mprj_la_data_in[117]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[117]/VPB ANTENNA_mprj_la_data_in[117]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[47] la_data_in[47] ANTENNA_mprj_la_data_in[47]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[47]/VPB ANTENNA_mprj_la_data_in[47]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[99] la_oen[99] ANTENNA_mprj_la_oen[99]/VGND VSUBS ANTENNA_mprj_la_oen[99]/VPB
+ ANTENNA_mprj_la_oen[99]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[27] wbs_adr_i[27] ANTENNA_mprj_wbs_adr_i[27]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[27]/VPB
+ ANTENNA_mprj_wbs_adr_i[27]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[23] io_in[23] ANTENNA_mprj_io_in[23]/VGND VSUBS ANTENNA_mprj_io_in[23]/VPB
+ ANTENNA_mprj_io_in[23]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[80] la_data_in[80] ANTENNA_mprj_la_data_in[80]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[80]/VPB ANTENNA_mprj_la_data_in[80]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[22] la_oen[22] ANTENNA_mprj_la_oen[22]/VGND VSUBS ANTENNA_mprj_la_oen[22]/VPB
+ ANTENNA_mprj_la_oen[22]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[63] la_data_in[63] ANTENNA_mprj_la_data_in[63]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[63]/VPB ANTENNA_mprj_la_data_in[63]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[46] la_data_in[46] ANTENNA_mprj_la_data_in[46]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[46]/VPB ANTENNA_mprj_la_data_in[46]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[116] la_data_in[116] ANTENNA_mprj_la_data_in[116]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[116]/VPB ANTENNA_mprj_la_data_in[116]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[29] la_data_in[29] ANTENNA_mprj_la_data_in[29]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[29]/VPB ANTENNA_mprj_la_data_in[29]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[26] wbs_adr_i[26] ANTENNA_mprj_wbs_adr_i[26]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[26]/VPB
+ ANTENNA_mprj_wbs_adr_i[26]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[22] io_in[22] ANTENNA_mprj_io_in[22]/VGND VSUBS ANTENNA_mprj_io_in[22]/VPB
+ ANTENNA_mprj_io_in[22]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[98] la_oen[98] ANTENNA_mprj_la_oen[98]/VGND VSUBS ANTENNA_mprj_la_oen[98]/VPB
+ ANTENNA_mprj_la_oen[98]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[21] la_oen[21] ANTENNA_mprj_la_oen[21]/VGND VSUBS ANTENNA_mprj_la_oen[21]/VPB
+ ANTENNA_mprj_la_oen[21]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[62] la_data_in[62] ANTENNA_mprj_la_data_in[62]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[62]/VPB ANTENNA_mprj_la_data_in[62]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wb_clk_i wb_clk_i ANTENNA_mprj_wb_clk_i/VGND VSUBS ANTENNA_mprj_wb_clk_i/VPB
+ ANTENNA_mprj_wb_clk_i/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[115] la_data_in[115] ANTENNA_mprj_la_data_in[115]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[115]/VPB ANTENNA_mprj_la_data_in[115]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[45] la_data_in[45] ANTENNA_mprj_la_data_in[45]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[45]/VPB ANTENNA_mprj_la_data_in[45]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[97] la_oen[97] ANTENNA_mprj_la_oen[97]/VGND VSUBS ANTENNA_mprj_la_oen[97]/VPB
+ ANTENNA_mprj_la_oen[97]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[28] la_data_in[28] ANTENNA_mprj_la_data_in[28]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[28]/VPB ANTENNA_mprj_la_data_in[28]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[25] wbs_adr_i[25] ANTENNA_mprj_wbs_adr_i[25]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[25]/VPB
+ ANTENNA_mprj_wbs_adr_i[25]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[21] io_in[21] ANTENNA_mprj_io_in[21]/VGND VSUBS ANTENNA_mprj_io_in[21]/VPB
+ ANTENNA_mprj_io_in[21]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[20] la_oen[20] ANTENNA_mprj_la_oen[20]/VGND VSUBS ANTENNA_mprj_la_oen[20]/VPB
+ ANTENNA_mprj_la_oen[20]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[61] la_data_in[61] ANTENNA_mprj_la_data_in[61]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[61]/VPB ANTENNA_mprj_la_data_in[61]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[44] la_data_in[44] ANTENNA_mprj_la_data_in[44]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[44]/VPB ANTENNA_mprj_la_data_in[44]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[114] la_data_in[114] ANTENNA_mprj_la_data_in[114]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[114]/VPB ANTENNA_mprj_la_data_in[114]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[27] la_data_in[27] ANTENNA_mprj_la_data_in[27]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[27]/VPB ANTENNA_mprj_la_data_in[27]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[24] wbs_adr_i[24] ANTENNA_mprj_wbs_adr_i[24]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[24]/VPB
+ ANTENNA_mprj_wbs_adr_i[24]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[96] la_oen[96] ANTENNA_mprj_la_oen[96]/VGND VSUBS ANTENNA_mprj_la_oen[96]/VPB
+ ANTENNA_mprj_la_oen[96]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[20] io_in[20] ANTENNA_mprj_io_in[20]/VGND VSUBS ANTENNA_mprj_io_in[20]/VPB
+ ANTENNA_mprj_io_in[20]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[79] la_oen[79] ANTENNA_mprj_la_oen[79]/VGND VSUBS ANTENNA_mprj_la_oen[79]/VPB
+ ANTENNA_mprj_la_oen[79]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[60] la_data_in[60] ANTENNA_mprj_la_data_in[60]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[60]/VPB ANTENNA_mprj_la_data_in[60]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[43] la_data_in[43] ANTENNA_mprj_la_data_in[43]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[43]/VPB ANTENNA_mprj_la_data_in[43]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_we_i wbs_we_i ANTENNA_mprj_wbs_we_i/VGND VSUBS ANTENNA_mprj_wbs_we_i/VPB
+ ANTENNA_mprj_wbs_we_i/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[113] la_data_in[113] ANTENNA_mprj_la_data_in[113]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[113]/VPB ANTENNA_mprj_la_data_in[113]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[95] la_oen[95] ANTENNA_mprj_la_oen[95]/VGND VSUBS ANTENNA_mprj_la_oen[95]/VPB
+ ANTENNA_mprj_la_oen[95]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[26] la_data_in[26] ANTENNA_mprj_la_data_in[26]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[26]/VPB ANTENNA_mprj_la_data_in[26]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[23] wbs_adr_i[23] ANTENNA_mprj_wbs_adr_i[23]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[23]/VPB
+ ANTENNA_mprj_wbs_adr_i[23]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[78] la_oen[78] ANTENNA_mprj_la_oen[78]/VGND VSUBS ANTENNA_mprj_la_oen[78]/VPB
+ ANTENNA_mprj_la_oen[78]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[19] wbs_dat_i[19] ANTENNA_mprj_wbs_dat_i[19]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[19]/VPB
+ ANTENNA_mprj_wbs_dat_i[19]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[112] la_data_in[112] ANTENNA_mprj_la_data_in[112]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[112]/VPB ANTENNA_mprj_la_data_in[112]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[42] la_data_in[42] ANTENNA_mprj_la_data_in[42]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[42]/VPB ANTENNA_mprj_la_data_in[42]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[25] la_data_in[25] ANTENNA_mprj_la_data_in[25]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[25]/VPB ANTENNA_mprj_la_data_in[25]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[94] la_oen[94] ANTENNA_mprj_la_oen[94]/VGND VSUBS ANTENNA_mprj_la_oen[94]/VPB
+ ANTENNA_mprj_la_oen[94]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[18] wbs_dat_i[18] ANTENNA_mprj_wbs_dat_i[18]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[18]/VPB
+ ANTENNA_mprj_wbs_dat_i[18]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[22] wbs_adr_i[22] ANTENNA_mprj_wbs_adr_i[22]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[22]/VPB
+ ANTENNA_mprj_wbs_adr_i[22]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[77] la_oen[77] ANTENNA_mprj_la_oen[77]/VGND VSUBS ANTENNA_mprj_la_oen[77]/VPB
+ ANTENNA_mprj_la_oen[77]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[41] la_data_in[41] ANTENNA_mprj_la_data_in[41]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[41]/VPB ANTENNA_mprj_la_data_in[41]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[111] la_data_in[111] ANTENNA_mprj_la_data_in[111]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[111]/VPB ANTENNA_mprj_la_data_in[111]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[24] la_data_in[24] ANTENNA_mprj_la_data_in[24]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[24]/VPB ANTENNA_mprj_la_data_in[24]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[21] wbs_adr_i[21] ANTENNA_mprj_wbs_adr_i[21]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[21]/VPB
+ ANTENNA_mprj_wbs_adr_i[21]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[119] la_oen[119] ANTENNA_mprj_la_oen[119]/VGND VSUBS ANTENNA_mprj_la_oen[119]/VPB
+ ANTENNA_mprj_la_oen[119]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[93] la_oen[93] ANTENNA_mprj_la_oen[93]/VGND VSUBS ANTENNA_mprj_la_oen[93]/VPB
+ ANTENNA_mprj_la_oen[93]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[76] la_oen[76] ANTENNA_mprj_la_oen[76]/VGND VSUBS ANTENNA_mprj_la_oen[76]/VPB
+ ANTENNA_mprj_la_oen[76]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[17] wbs_dat_i[17] ANTENNA_mprj_wbs_dat_i[17]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[17]/VPB
+ ANTENNA_mprj_wbs_dat_i[17]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[59] la_oen[59] ANTENNA_mprj_la_oen[59]/VGND VSUBS ANTENNA_mprj_la_oen[59]/VPB
+ ANTENNA_mprj_la_oen[59]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[110] la_data_in[110] ANTENNA_mprj_la_data_in[110]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[110]/VPB ANTENNA_mprj_la_data_in[110]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[40] la_data_in[40] ANTENNA_mprj_la_data_in[40]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[40]/VPB ANTENNA_mprj_la_data_in[40]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[23] la_data_in[23] ANTENNA_mprj_la_data_in[23]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[23]/VPB ANTENNA_mprj_la_data_in[23]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[118] la_oen[118] ANTENNA_mprj_la_oen[118]/VGND VSUBS ANTENNA_mprj_la_oen[118]/VPB
+ ANTENNA_mprj_la_oen[118]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[92] la_oen[92] ANTENNA_mprj_la_oen[92]/VGND VSUBS ANTENNA_mprj_la_oen[92]/VPB
+ ANTENNA_mprj_la_oen[92]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[16] wbs_dat_i[16] ANTENNA_mprj_wbs_dat_i[16]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[16]/VPB
+ ANTENNA_mprj_wbs_dat_i[16]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[20] wbs_adr_i[20] ANTENNA_mprj_wbs_adr_i[20]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[20]/VPB
+ ANTENNA_mprj_wbs_adr_i[20]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[75] la_oen[75] ANTENNA_mprj_la_oen[75]/VGND VSUBS ANTENNA_mprj_la_oen[75]/VPB
+ ANTENNA_mprj_la_oen[75]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[58] la_oen[58] ANTENNA_mprj_la_oen[58]/VGND VSUBS ANTENNA_mprj_la_oen[58]/VPB
+ ANTENNA_mprj_la_oen[58]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[99] la_data_in[99] ANTENNA_mprj_la_data_in[99]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[99]/VPB ANTENNA_mprj_la_data_in[99]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[22] la_data_in[22] ANTENNA_mprj_la_data_in[22]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[22]/VPB ANTENNA_mprj_la_data_in[22]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[117] la_oen[117] ANTENNA_mprj_la_oen[117]/VGND VSUBS ANTENNA_mprj_la_oen[117]/VPB
+ ANTENNA_mprj_la_oen[117]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[91] la_oen[91] ANTENNA_mprj_la_oen[91]/VGND VSUBS ANTENNA_mprj_la_oen[91]/VPB
+ ANTENNA_mprj_la_oen[91]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[74] la_oen[74] ANTENNA_mprj_la_oen[74]/VGND VSUBS ANTENNA_mprj_la_oen[74]/VPB
+ ANTENNA_mprj_la_oen[74]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[15] wbs_dat_i[15] ANTENNA_mprj_wbs_dat_i[15]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[15]/VPB
+ ANTENNA_mprj_wbs_dat_i[15]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[57] la_oen[57] ANTENNA_mprj_la_oen[57]/VGND VSUBS ANTENNA_mprj_la_oen[57]/VPB
+ ANTENNA_mprj_la_oen[57]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[98] la_data_in[98] ANTENNA_mprj_la_data_in[98]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[98]/VPB ANTENNA_mprj_la_data_in[98]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[21] la_data_in[21] ANTENNA_mprj_la_data_in[21]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[21]/VPB ANTENNA_mprj_la_data_in[21]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[9] la_data_in[9] ANTENNA_mprj_la_data_in[9]/VGND VSUBS ANTENNA_mprj_la_data_in[9]/VPB
+ ANTENNA_mprj_la_data_in[9]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[116] la_oen[116] ANTENNA_mprj_la_oen[116]/VGND VSUBS ANTENNA_mprj_la_oen[116]/VPB
+ ANTENNA_mprj_la_oen[116]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[90] la_oen[90] ANTENNA_mprj_la_oen[90]/VGND VSUBS ANTENNA_mprj_la_oen[90]/VPB
+ ANTENNA_mprj_la_oen[90]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[14] wbs_dat_i[14] ANTENNA_mprj_wbs_dat_i[14]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[14]/VPB
+ ANTENNA_mprj_wbs_dat_i[14]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[31] wbs_dat_i[31] ANTENNA_mprj_wbs_dat_i[31]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[31]/VPB
+ ANTENNA_mprj_wbs_dat_i[31]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[73] la_oen[73] ANTENNA_mprj_la_oen[73]/VGND VSUBS ANTENNA_mprj_la_oen[73]/VPB
+ ANTENNA_mprj_la_oen[73]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[56] la_oen[56] ANTENNA_mprj_la_oen[56]/VGND VSUBS ANTENNA_mprj_la_oen[56]/VPB
+ ANTENNA_mprj_la_oen[56]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[39] la_oen[39] ANTENNA_mprj_la_oen[39]/VGND VSUBS ANTENNA_mprj_la_oen[39]/VPB
+ ANTENNA_mprj_la_oen[39]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[97] la_data_in[97] ANTENNA_mprj_la_data_in[97]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[97]/VPB ANTENNA_mprj_la_data_in[97]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[20] la_data_in[20] ANTENNA_mprj_la_data_in[20]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[20]/VPB ANTENNA_mprj_la_data_in[20]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[30] wbs_dat_i[30] ANTENNA_mprj_wbs_dat_i[30]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[30]/VPB
+ ANTENNA_mprj_wbs_dat_i[30]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[8] la_data_in[8] ANTENNA_mprj_la_data_in[8]/VGND VSUBS ANTENNA_mprj_la_data_in[8]/VPB
+ ANTENNA_mprj_la_data_in[8]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[115] la_oen[115] ANTENNA_mprj_la_oen[115]/VGND VSUBS ANTENNA_mprj_la_oen[115]/VPB
+ ANTENNA_mprj_la_oen[115]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[72] la_oen[72] ANTENNA_mprj_la_oen[72]/VGND VSUBS ANTENNA_mprj_la_oen[72]/VPB
+ ANTENNA_mprj_la_oen[72]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[13] wbs_dat_i[13] ANTENNA_mprj_wbs_dat_i[13]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[13]/VPB
+ ANTENNA_mprj_wbs_dat_i[13]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[55] la_oen[55] ANTENNA_mprj_la_oen[55]/VGND VSUBS ANTENNA_mprj_la_oen[55]/VPB
+ ANTENNA_mprj_la_oen[55]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[96] la_data_in[96] ANTENNA_mprj_la_data_in[96]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[96]/VPB ANTENNA_mprj_la_data_in[96]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[38] la_oen[38] ANTENNA_mprj_la_oen[38]/VGND VSUBS ANTENNA_mprj_la_oen[38]/VPB
+ ANTENNA_mprj_la_oen[38]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[7] la_data_in[7] ANTENNA_mprj_la_data_in[7]/VGND VSUBS ANTENNA_mprj_la_data_in[7]/VPB
+ ANTENNA_mprj_la_data_in[7]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[79] la_data_in[79] ANTENNA_mprj_la_data_in[79]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[79]/VPB ANTENNA_mprj_la_data_in[79]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[12] wbs_dat_i[12] ANTENNA_mprj_wbs_dat_i[12]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[12]/VPB
+ ANTENNA_mprj_wbs_dat_i[12]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[114] la_oen[114] ANTENNA_mprj_la_oen[114]/VGND VSUBS ANTENNA_mprj_la_oen[114]/VPB
+ ANTENNA_mprj_la_oen[114]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[71] la_oen[71] ANTENNA_mprj_la_oen[71]/VGND VSUBS ANTENNA_mprj_la_oen[71]/VPB
+ ANTENNA_mprj_la_oen[71]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[54] la_oen[54] ANTENNA_mprj_la_oen[54]/VGND VSUBS ANTENNA_mprj_la_oen[54]/VPB
+ ANTENNA_mprj_la_oen[54]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[37] la_oen[37] ANTENNA_mprj_la_oen[37]/VGND VSUBS ANTENNA_mprj_la_oen[37]/VPB
+ ANTENNA_mprj_la_oen[37]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[95] la_data_in[95] ANTENNA_mprj_la_data_in[95]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[95]/VPB ANTENNA_mprj_la_data_in[95]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[78] la_data_in[78] ANTENNA_mprj_la_data_in[78]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[78]/VPB ANTENNA_mprj_la_data_in[78]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[6] la_data_in[6] ANTENNA_mprj_la_data_in[6]/VGND VSUBS ANTENNA_mprj_la_data_in[6]/VPB
+ ANTENNA_mprj_la_data_in[6]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[113] la_oen[113] ANTENNA_mprj_la_oen[113]/VGND VSUBS ANTENNA_mprj_la_oen[113]/VPB
+ ANTENNA_mprj_la_oen[113]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[70] la_oen[70] ANTENNA_mprj_la_oen[70]/VGND VSUBS ANTENNA_mprj_la_oen[70]/VPB
+ ANTENNA_mprj_la_oen[70]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[11] wbs_dat_i[11] ANTENNA_mprj_wbs_dat_i[11]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[11]/VPB
+ ANTENNA_mprj_wbs_dat_i[11]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[9] io_in[9] ANTENNA_mprj_io_in[9]/VGND VSUBS ANTENNA_mprj_io_in[9]/VPB
+ ANTENNA_mprj_io_in[9]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[53] la_oen[53] ANTENNA_mprj_la_oen[53]/VGND VSUBS ANTENNA_mprj_la_oen[53]/VPB
+ ANTENNA_mprj_la_oen[53]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[94] la_data_in[94] ANTENNA_mprj_la_data_in[94]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[94]/VPB ANTENNA_mprj_la_data_in[94]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[36] la_oen[36] ANTENNA_mprj_la_oen[36]/VGND VSUBS ANTENNA_mprj_la_oen[36]/VPB
+ ANTENNA_mprj_la_oen[36]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[37] io_in[37] ANTENNA_mprj_io_in[37]/VGND VSUBS ANTENNA_mprj_io_in[37]/VPB
+ ANTENNA_mprj_io_in[37]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[5] la_data_in[5] ANTENNA_mprj_la_data_in[5]/VGND VSUBS ANTENNA_mprj_la_data_in[5]/VPB
+ ANTENNA_mprj_la_data_in[5]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[77] la_data_in[77] ANTENNA_mprj_la_data_in[77]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[77]/VPB ANTENNA_mprj_la_data_in[77]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[19] la_oen[19] ANTENNA_mprj_la_oen[19]/VGND VSUBS ANTENNA_mprj_la_oen[19]/VPB
+ ANTENNA_mprj_la_oen[19]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[10] wbs_dat_i[10] ANTENNA_mprj_wbs_dat_i[10]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[10]/VPB
+ ANTENNA_mprj_wbs_dat_i[10]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[112] la_oen[112] ANTENNA_mprj_la_oen[112]/VGND VSUBS ANTENNA_mprj_la_oen[112]/VPB
+ ANTENNA_mprj_la_oen[112]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[8] io_in[8] ANTENNA_mprj_io_in[8]/VGND VSUBS ANTENNA_mprj_io_in[8]/VPB
+ ANTENNA_mprj_io_in[8]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[52] la_oen[52] ANTENNA_mprj_la_oen[52]/VGND VSUBS ANTENNA_mprj_la_oen[52]/VPB
+ ANTENNA_mprj_la_oen[52]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[35] la_oen[35] ANTENNA_mprj_la_oen[35]/VGND VSUBS ANTENNA_mprj_la_oen[35]/VPB
+ ANTENNA_mprj_la_oen[35]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[19] io_in[19] ANTENNA_mprj_io_in[19]/VGND VSUBS ANTENNA_mprj_io_in[19]/VPB
+ ANTENNA_mprj_io_in[19]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[36] io_in[36] ANTENNA_mprj_io_in[36]/VGND VSUBS ANTENNA_mprj_io_in[36]/VPB
+ ANTENNA_mprj_io_in[36]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[93] la_data_in[93] ANTENNA_mprj_la_data_in[93]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[93]/VPB ANTENNA_mprj_la_data_in[93]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[76] la_data_in[76] ANTENNA_mprj_la_data_in[76]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[76]/VPB ANTENNA_mprj_la_data_in[76]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[18] la_oen[18] ANTENNA_mprj_la_oen[18]/VGND VSUBS ANTENNA_mprj_la_oen[18]/VPB
+ ANTENNA_mprj_la_oen[18]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[4] la_data_in[4] ANTENNA_mprj_la_data_in[4]/VGND VSUBS ANTENNA_mprj_la_data_in[4]/VPB
+ ANTENNA_mprj_la_data_in[4]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[111] la_oen[111] ANTENNA_mprj_la_oen[111]/VGND VSUBS ANTENNA_mprj_la_oen[111]/VPB
+ ANTENNA_mprj_la_oen[111]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[59] la_data_in[59] ANTENNA_mprj_la_data_in[59]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[59]/VPB ANTENNA_mprj_la_data_in[59]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[7] io_in[7] ANTENNA_mprj_io_in[7]/VGND VSUBS ANTENNA_mprj_io_in[7]/VPB
+ ANTENNA_mprj_io_in[7]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[51] la_oen[51] ANTENNA_mprj_la_oen[51]/VGND VSUBS ANTENNA_mprj_la_oen[51]/VPB
+ ANTENNA_mprj_la_oen[51]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[35] io_in[35] ANTENNA_mprj_io_in[35]/VGND VSUBS ANTENNA_mprj_io_in[35]/VPB
+ ANTENNA_mprj_io_in[35]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[92] la_data_in[92] ANTENNA_mprj_la_data_in[92]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[92]/VPB ANTENNA_mprj_la_data_in[92]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[34] la_oen[34] ANTENNA_mprj_la_oen[34]/VGND VSUBS ANTENNA_mprj_la_oen[34]/VPB
+ ANTENNA_mprj_la_oen[34]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[3] la_data_in[3] ANTENNA_mprj_la_data_in[3]/VGND VSUBS ANTENNA_mprj_la_data_in[3]/VPB
+ ANTENNA_mprj_la_data_in[3]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[18] io_in[18] ANTENNA_mprj_io_in[18]/VGND VSUBS ANTENNA_mprj_io_in[18]/VPB
+ ANTENNA_mprj_io_in[18]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[75] la_data_in[75] ANTENNA_mprj_la_data_in[75]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[75]/VPB ANTENNA_mprj_la_data_in[75]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[17] la_oen[17] ANTENNA_mprj_la_oen[17]/VGND VSUBS ANTENNA_mprj_la_oen[17]/VPB
+ ANTENNA_mprj_la_oen[17]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[110] la_oen[110] ANTENNA_mprj_la_oen[110]/VGND VSUBS ANTENNA_mprj_la_oen[110]/VPB
+ ANTENNA_mprj_la_oen[110]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[58] la_data_in[58] ANTENNA_mprj_la_data_in[58]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[58]/VPB ANTENNA_mprj_la_data_in[58]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[6] io_in[6] ANTENNA_mprj_io_in[6]/VGND VSUBS ANTENNA_mprj_io_in[6]/VPB
+ ANTENNA_mprj_io_in[6]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[50] la_oen[50] ANTENNA_mprj_la_oen[50]/VGND VSUBS ANTENNA_mprj_la_oen[50]/VPB
+ ANTENNA_mprj_la_oen[50]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[33] la_oen[33] ANTENNA_mprj_la_oen[33]/VGND VSUBS ANTENNA_mprj_la_oen[33]/VPB
+ ANTENNA_mprj_la_oen[33]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_stb_i wbs_stb_i ANTENNA_mprj_wbs_stb_i/VGND VSUBS ANTENNA_mprj_wbs_stb_i/VPB
+ ANTENNA_mprj_wbs_stb_i/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[17] io_in[17] ANTENNA_mprj_io_in[17]/VGND VSUBS ANTENNA_mprj_io_in[17]/VPB
+ ANTENNA_mprj_io_in[17]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[34] io_in[34] ANTENNA_mprj_io_in[34]/VGND VSUBS ANTENNA_mprj_io_in[34]/VPB
+ ANTENNA_mprj_io_in[34]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[91] la_data_in[91] ANTENNA_mprj_la_data_in[91]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[91]/VPB ANTENNA_mprj_la_data_in[91]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[74] la_data_in[74] ANTENNA_mprj_la_data_in[74]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[74]/VPB ANTENNA_mprj_la_data_in[74]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[16] la_oen[16] ANTENNA_mprj_la_oen[16]/VGND VSUBS ANTENNA_mprj_la_oen[16]/VPB
+ ANTENNA_mprj_la_oen[16]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[2] la_data_in[2] ANTENNA_mprj_la_data_in[2]/VGND VSUBS ANTENNA_mprj_la_data_in[2]/VPB
+ ANTENNA_mprj_la_data_in[2]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[57] la_data_in[57] ANTENNA_mprj_la_data_in[57]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[57]/VPB ANTENNA_mprj_la_data_in[57]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[127] la_data_in[127] ANTENNA_mprj_la_oen[127]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[127]/VPB ANTENNA_mprj_la_data_in[127]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[5] io_in[5] ANTENNA_mprj_io_in[5]/VGND VSUBS ANTENNA_mprj_io_in[5]/VPB
+ ANTENNA_mprj_io_in[5]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[33] io_in[33] ANTENNA_mprj_io_in[33]/VGND VSUBS ANTENNA_mprj_io_in[33]/VPB
+ ANTENNA_mprj_io_in[33]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[90] la_data_in[90] ANTENNA_mprj_la_data_in[90]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[90]/VPB ANTENNA_mprj_la_data_in[90]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[32] la_oen[32] ANTENNA_mprj_la_oen[32]/VGND VSUBS ANTENNA_mprj_la_oen[32]/VPB
+ ANTENNA_mprj_la_oen[32]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[16] io_in[16] ANTENNA_mprj_io_in[16]/VGND VSUBS ANTENNA_mprj_io_in[16]/VPB
+ ANTENNA_mprj_io_in[16]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[73] la_data_in[73] ANTENNA_mprj_la_data_in[73]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[73]/VPB ANTENNA_mprj_la_data_in[73]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[15] la_oen[15] ANTENNA_mprj_la_oen[15]/VGND VSUBS ANTENNA_mprj_la_oen[15]/VPB
+ ANTENNA_mprj_la_oen[15]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[1] la_data_in[1] ANTENNA_mprj_la_data_in[1]/VGND VSUBS ANTENNA_mprj_la_data_in[1]/VPB
+ ANTENNA_mprj_la_data_in[1]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[126] la_data_in[126] ANTENNA_mprj_la_data_in[126]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[126]/VPB ANTENNA_mprj_la_data_in[126]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[56] la_data_in[56] ANTENNA_mprj_la_data_in[56]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[56]/VPB ANTENNA_mprj_la_data_in[56]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[39] la_data_in[39] ANTENNA_mprj_la_data_in[39]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[39]/VPB ANTENNA_mprj_la_data_in[39]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[4] io_in[4] ANTENNA_mprj_io_in[4]/VGND VSUBS ANTENNA_mprj_io_in[4]/VPB
+ ANTENNA_mprj_io_in[4]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[109] la_data_in[109] ANTENNA_mprj_la_data_in[109]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[109]/VPB ANTENNA_mprj_la_data_in[109]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[19] wbs_adr_i[19] ANTENNA_mprj_wbs_adr_i[19]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[19]/VPB
+ ANTENNA_mprj_wbs_adr_i[19]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[15] io_in[15] ANTENNA_mprj_io_in[15]/VGND VSUBS ANTENNA_mprj_io_in[15]/VPB
+ ANTENNA_mprj_io_in[15]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[32] io_in[32] ANTENNA_mprj_io_in[32]/VGND VSUBS ANTENNA_mprj_io_in[32]/VPB
+ ANTENNA_mprj_io_in[32]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[31] la_oen[31] ANTENNA_mprj_la_oen[31]/VGND VSUBS ANTENNA_mprj_la_oen[31]/VPB
+ ANTENNA_mprj_la_oen[31]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[14] la_oen[14] ANTENNA_mprj_la_oen[14]/VGND VSUBS ANTENNA_mprj_la_oen[14]/VPB
+ ANTENNA_mprj_la_oen[14]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_cyc_i wbs_cyc_i ANTENNA_mprj_wbs_cyc_i/VGND VSUBS ANTENNA_mprj_wbs_cyc_i/VPB
+ ANTENNA_mprj_wbs_cyc_i/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[0] la_data_in[0] ANTENNA_mprj_la_data_in[0]/VGND VSUBS ANTENNA_mprj_la_data_in[0]/VPB
+ ANTENNA_mprj_la_data_in[0]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[72] la_data_in[72] ANTENNA_mprj_la_data_in[72]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[72]/VPB ANTENNA_mprj_la_data_in[72]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[55] la_data_in[55] ANTENNA_mprj_la_data_in[55]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[55]/VPB ANTENNA_mprj_la_data_in[55]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[125] la_data_in[125] ANTENNA_mprj_la_data_in[125]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[125]/VPB ANTENNA_mprj_la_data_in[125]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[108] la_data_in[108] ANTENNA_mprj_la_data_in[108]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[108]/VPB ANTENNA_mprj_la_data_in[108]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[38] la_data_in[38] ANTENNA_mprj_la_data_in[38]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[38]/VPB ANTENNA_mprj_la_data_in[38]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[31] io_in[31] ANTENNA_mprj_io_in[31]/VGND VSUBS ANTENNA_mprj_io_in[31]/VPB
+ ANTENNA_mprj_io_in[31]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[3] io_in[3] ANTENNA_mprj_io_in[3]/VGND VSUBS ANTENNA_mprj_io_in[3]/VPB
+ ANTENNA_mprj_io_in[3]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[30] la_oen[30] ANTENNA_mprj_la_oen[30]/VGND VSUBS ANTENNA_mprj_la_oen[30]/VPB
+ ANTENNA_mprj_la_oen[30]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[18] wbs_adr_i[18] ANTENNA_mprj_wbs_adr_i[18]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[18]/VPB
+ ANTENNA_mprj_wbs_adr_i[18]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[14] io_in[14] ANTENNA_mprj_io_in[14]/VGND VSUBS ANTENNA_mprj_io_in[14]/VPB
+ ANTENNA_mprj_io_in[14]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[71] la_data_in[71] ANTENNA_mprj_la_data_in[71]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[71]/VPB ANTENNA_mprj_la_data_in[71]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[13] la_oen[13] ANTENNA_mprj_la_oen[13]/VGND VSUBS ANTENNA_mprj_la_oen[13]/VPB
+ ANTENNA_mprj_la_oen[13]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[9] wbs_adr_i[9] ANTENNA_mprj_wbs_adr_i[9]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[9]/VPB
+ ANTENNA_mprj_wbs_adr_i[9]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[124] la_data_in[124] ANTENNA_mprj_la_data_in[124]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[124]/VPB ANTENNA_mprj_la_data_in[124]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[54] la_data_in[54] ANTENNA_mprj_la_data_in[54]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[54]/VPB ANTENNA_mprj_la_data_in[54]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[37] la_data_in[37] ANTENNA_mprj_la_data_in[37]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[37]/VPB ANTENNA_mprj_la_data_in[37]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[2] io_in[2] ANTENNA_mprj_io_in[2]/VGND VSUBS ANTENNA_mprj_io_in[2]/VPB
+ ANTENNA_mprj_io_in[2]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[107] la_data_in[107] ANTENNA_mprj_la_data_in[107]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[107]/VPB ANTENNA_mprj_la_data_in[107]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[17] wbs_adr_i[17] ANTENNA_mprj_wbs_adr_i[17]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[17]/VPB
+ ANTENNA_mprj_wbs_adr_i[17]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[30] io_in[30] ANTENNA_mprj_io_in[30]/VGND VSUBS ANTENNA_mprj_io_in[30]/VPB
+ ANTENNA_mprj_io_in[30]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[89] la_oen[89] ANTENNA_mprj_la_oen[89]/VGND VSUBS ANTENNA_mprj_la_oen[89]/VPB
+ ANTENNA_mprj_la_oen[89]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[12] la_oen[12] ANTENNA_mprj_la_oen[12]/VGND VSUBS ANTENNA_mprj_la_oen[12]/VPB
+ ANTENNA_mprj_la_oen[12]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[9] wbs_dat_i[9] ANTENNA_mprj_wbs_dat_i[9]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[9]/VPB
+ ANTENNA_mprj_wbs_dat_i[9]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[13] io_in[13] ANTENNA_mprj_io_in[13]/VGND VSUBS ANTENNA_mprj_io_in[13]/VPB
+ ANTENNA_mprj_io_in[13]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[70] la_data_in[70] ANTENNA_mprj_la_data_in[70]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[70]/VPB ANTENNA_mprj_la_data_in[70]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[53] la_data_in[53] ANTENNA_mprj_la_data_in[53]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[53]/VPB ANTENNA_mprj_la_data_in[53]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[8] wbs_adr_i[8] ANTENNA_mprj_wbs_adr_i[8]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[8]/VPB
+ ANTENNA_mprj_wbs_adr_i[8]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[123] la_data_in[123] ANTENNA_mprj_la_data_in[123]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[123]/VPB ANTENNA_mprj_la_data_in[123]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[36] la_data_in[36] ANTENNA_mprj_la_data_in[36]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[36]/VPB ANTENNA_mprj_la_data_in[36]/VPWR sky130_fd_sc_hd__diode_2
Xmprj io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16]
+ io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24]
+ io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32]
+ io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20]
+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28]
+ io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35]
+ io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2]
+ io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0]
+ la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oen[0] la_oen[100] la_oen[101]
+ la_oen[102] la_oen[103] la_oen[104] la_oen[105] la_oen[106] la_oen[107] la_oen[108]
+ la_oen[109] la_oen[10] la_oen[110] la_oen[111] la_oen[112] la_oen[113] la_oen[114]
+ la_oen[115] la_oen[116] la_oen[117] la_oen[118] la_oen[119] la_oen[11] la_oen[120]
+ la_oen[121] la_oen[122] la_oen[123] la_oen[124] la_oen[125] la_oen[126] la_oen[127]
+ la_oen[12] la_oen[13] la_oen[14] la_oen[15] la_oen[16] la_oen[17] la_oen[18] la_oen[19]
+ la_oen[1] la_oen[20] la_oen[21] la_oen[22] la_oen[23] la_oen[24] la_oen[25] la_oen[26]
+ la_oen[27] la_oen[28] la_oen[29] la_oen[2] la_oen[30] la_oen[31] la_oen[32] la_oen[33]
+ la_oen[34] la_oen[35] la_oen[36] la_oen[37] la_oen[38] la_oen[39] la_oen[3] la_oen[40]
+ la_oen[41] la_oen[42] la_oen[43] la_oen[44] la_oen[45] la_oen[46] la_oen[47] la_oen[48]
+ la_oen[49] la_oen[4] la_oen[50] la_oen[51] la_oen[52] la_oen[53] la_oen[54] la_oen[55]
+ la_oen[56] la_oen[57] la_oen[58] la_oen[59] la_oen[5] la_oen[60] la_oen[61] la_oen[62]
+ la_oen[63] la_oen[64] la_oen[65] la_oen[66] la_oen[67] la_oen[68] la_oen[69] la_oen[6]
+ la_oen[70] la_oen[71] la_oen[72] la_oen[73] la_oen[74] la_oen[75] la_oen[76] la_oen[77]
+ la_oen[78] la_oen[79] la_oen[7] la_oen[80] la_oen[81] la_oen[82] la_oen[83] la_oen[84]
+ la_oen[85] la_oen[86] la_oen[87] la_oen[88] la_oen[89] la_oen[8] la_oen[90] la_oen[91]
+ la_oen[92] la_oen[93] la_oen[94] la_oen[95] la_oen[96] la_oen[97] la_oen[98] la_oen[99]
+ la_oen[9] wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i mprj/VPWR
+ mprj/VGND accelerator_top
XANTENNA_mprj_io_in[1] io_in[1] ANTENNA_mprj_io_in[1]/VGND VSUBS ANTENNA_mprj_io_in[1]/VPB
+ ANTENNA_mprj_io_in[1]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[106] la_data_in[106] ANTENNA_mprj_la_data_in[106]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[106]/VPB ANTENNA_mprj_la_data_in[106]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[88] la_oen[88] ANTENNA_mprj_la_oen[88]/VGND VSUBS ANTENNA_mprj_la_oen[88]/VPB
+ ANTENNA_mprj_la_oen[88]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[19] la_data_in[19] ANTENNA_mprj_la_data_in[19]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[19]/VPB ANTENNA_mprj_la_data_in[19]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[16] wbs_adr_i[16] ANTENNA_mprj_wbs_adr_i[16]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[16]/VPB
+ ANTENNA_mprj_wbs_adr_i[16]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[29] wbs_dat_i[29] ANTENNA_mprj_wbs_dat_i[29]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[29]/VPB
+ ANTENNA_mprj_wbs_dat_i[29]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[12] io_in[12] ANTENNA_mprj_io_in[12]/VGND VSUBS ANTENNA_mprj_io_in[12]/VPB
+ ANTENNA_mprj_io_in[12]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[11] la_oen[11] ANTENNA_mprj_la_oen[11]/VGND VSUBS ANTENNA_mprj_la_oen[11]/VPB
+ ANTENNA_mprj_la_oen[11]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[7] wbs_adr_i[7] ANTENNA_mprj_wbs_adr_i[7]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[7]/VPB
+ ANTENNA_mprj_wbs_adr_i[7]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[8] wbs_dat_i[8] ANTENNA_mprj_wbs_dat_i[8]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[8]/VPB
+ ANTENNA_mprj_wbs_dat_i[8]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[122] la_data_in[122] ANTENNA_mprj_la_data_in[122]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[122]/VPB ANTENNA_mprj_la_data_in[122]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[52] la_data_in[52] ANTENNA_mprj_la_data_in[52]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[52]/VPB ANTENNA_mprj_la_data_in[52]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[0] io_in[0] ANTENNA_mprj_io_in[0]/VGND VSUBS ANTENNA_mprj_io_in[0]/VPB
+ ANTENNA_mprj_io_in[0]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[105] la_data_in[105] ANTENNA_mprj_la_data_in[105]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[105]/VPB ANTENNA_mprj_la_data_in[105]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[35] la_data_in[35] ANTENNA_mprj_la_data_in[35]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[35]/VPB ANTENNA_mprj_la_data_in[35]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[18] la_data_in[18] ANTENNA_mprj_la_data_in[18]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[18]/VPB ANTENNA_mprj_la_data_in[18]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[28] wbs_dat_i[28] ANTENNA_mprj_wbs_dat_i[28]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[28]/VPB
+ ANTENNA_mprj_wbs_dat_i[28]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[87] la_oen[87] ANTENNA_mprj_la_oen[87]/VGND VSUBS ANTENNA_mprj_la_oen[87]/VPB
+ ANTENNA_mprj_la_oen[87]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[10] la_oen[10] ANTENNA_mprj_la_oen[10]/VGND VSUBS ANTENNA_mprj_la_oen[10]/VPB
+ ANTENNA_mprj_la_oen[10]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[15] wbs_adr_i[15] ANTENNA_mprj_wbs_adr_i[15]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[15]/VPB
+ ANTENNA_mprj_wbs_adr_i[15]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[11] io_in[11] ANTENNA_mprj_io_in[11]/VGND VSUBS ANTENNA_mprj_io_in[11]/VPB
+ ANTENNA_mprj_io_in[11]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[51] la_data_in[51] ANTENNA_mprj_la_data_in[51]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[51]/VPB ANTENNA_mprj_la_data_in[51]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[6] wbs_adr_i[6] ANTENNA_mprj_wbs_adr_i[6]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[6]/VPB
+ ANTENNA_mprj_wbs_adr_i[6]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[7] wbs_dat_i[7] ANTENNA_mprj_wbs_dat_i[7]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[7]/VPB
+ ANTENNA_mprj_wbs_dat_i[7]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[121] la_data_in[121] ANTENNA_mprj_la_data_in[121]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[121]/VPB ANTENNA_mprj_la_data_in[121]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[34] la_data_in[34] ANTENNA_mprj_la_data_in[34]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[34]/VPB ANTENNA_mprj_la_data_in[34]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[31] wbs_adr_i[31] ANTENNA_mprj_wbs_adr_i[31]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[31]/VPB
+ ANTENNA_mprj_wbs_adr_i[31]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[104] la_data_in[104] ANTENNA_mprj_la_data_in[104]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[104]/VPB ANTENNA_mprj_la_data_in[104]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[17] la_data_in[17] ANTENNA_mprj_la_data_in[17]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[17]/VPB ANTENNA_mprj_la_data_in[17]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[14] wbs_adr_i[14] ANTENNA_mprj_wbs_adr_i[14]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[14]/VPB
+ ANTENNA_mprj_wbs_adr_i[14]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[27] wbs_dat_i[27] ANTENNA_mprj_wbs_dat_i[27]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[27]/VPB
+ ANTENNA_mprj_wbs_dat_i[27]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[9] la_oen[9] ANTENNA_mprj_la_oen[9]/VGND VSUBS ANTENNA_mprj_la_oen[9]/VPB
+ ANTENNA_mprj_la_oen[9]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_io_in[10] io_in[10] ANTENNA_mprj_io_in[10]/VGND VSUBS ANTENNA_mprj_io_in[10]/VPB
+ ANTENNA_mprj_io_in[10]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[86] la_oen[86] ANTENNA_mprj_la_oen[86]/VGND VSUBS ANTENNA_mprj_la_oen[86]/VPB
+ ANTENNA_mprj_la_oen[86]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[69] la_oen[69] ANTENNA_mprj_la_oen[69]/VGND VSUBS ANTENNA_mprj_la_oen[69]/VPB
+ ANTENNA_mprj_la_oen[69]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[5] wbs_adr_i[5] ANTENNA_mprj_wbs_adr_i[5]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[5]/VPB
+ ANTENNA_mprj_wbs_adr_i[5]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[6] wbs_dat_i[6] ANTENNA_mprj_wbs_dat_i[6]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[6]/VPB
+ ANTENNA_mprj_wbs_dat_i[6]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[50] la_data_in[50] ANTENNA_mprj_la_data_in[50]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[50]/VPB ANTENNA_mprj_la_data_in[50]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[120] la_data_in[120] ANTENNA_mprj_la_data_in[120]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[120]/VPB ANTENNA_mprj_la_data_in[120]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[103] la_data_in[103] ANTENNA_mprj_la_data_in[103]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[103]/VPB ANTENNA_mprj_la_data_in[103]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[33] la_data_in[33] ANTENNA_mprj_la_data_in[33]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[33]/VPB ANTENNA_mprj_la_data_in[33]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[16] la_data_in[16] ANTENNA_mprj_la_data_in[16]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[16]/VPB ANTENNA_mprj_la_data_in[16]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[30] wbs_adr_i[30] ANTENNA_mprj_wbs_adr_i[30]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[30]/VPB
+ ANTENNA_mprj_wbs_adr_i[30]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[85] la_oen[85] ANTENNA_mprj_la_oen[85]/VGND VSUBS ANTENNA_mprj_la_oen[85]/VPB
+ ANTENNA_mprj_la_oen[85]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[13] wbs_adr_i[13] ANTENNA_mprj_wbs_adr_i[13]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[13]/VPB
+ ANTENNA_mprj_wbs_adr_i[13]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[26] wbs_dat_i[26] ANTENNA_mprj_wbs_dat_i[26]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[26]/VPB
+ ANTENNA_mprj_wbs_dat_i[26]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[8] la_oen[8] ANTENNA_mprj_la_oen[8]/VGND VSUBS ANTENNA_mprj_la_oen[8]/VPB
+ ANTENNA_mprj_la_oen[8]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[68] la_oen[68] ANTENNA_mprj_la_oen[68]/VGND VSUBS ANTENNA_mprj_la_oen[68]/VPB
+ ANTENNA_mprj_la_oen[68]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[4] wbs_adr_i[4] ANTENNA_mprj_wbs_adr_i[4]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[4]/VPB
+ ANTENNA_mprj_wbs_adr_i[4]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[5] wbs_dat_i[5] ANTENNA_mprj_wbs_dat_i[5]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[5]/VPB
+ ANTENNA_mprj_wbs_dat_i[5]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[32] la_data_in[32] ANTENNA_mprj_la_data_in[32]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[32]/VPB ANTENNA_mprj_la_data_in[32]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[127] la_oen[127] ANTENNA_mprj_la_oen[127]/VGND VSUBS ANTENNA_mprj_la_oen[127]/VPB
+ ANTENNA_mprj_la_oen[127]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[102] la_data_in[102] ANTENNA_mprj_la_data_in[102]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[102]/VPB ANTENNA_mprj_la_data_in[102]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[15] la_data_in[15] ANTENNA_mprj_la_data_in[15]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[15]/VPB ANTENNA_mprj_la_data_in[15]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[12] wbs_adr_i[12] ANTENNA_mprj_wbs_adr_i[12]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[12]/VPB
+ ANTENNA_mprj_wbs_adr_i[12]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[25] wbs_dat_i[25] ANTENNA_mprj_wbs_dat_i[25]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[25]/VPB
+ ANTENNA_mprj_wbs_dat_i[25]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[7] la_oen[7] ANTENNA_mprj_la_oen[7]/VGND VSUBS ANTENNA_mprj_la_oen[7]/VPB
+ ANTENNA_mprj_la_oen[7]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[84] la_oen[84] ANTENNA_mprj_la_oen[84]/VGND VSUBS ANTENNA_mprj_la_oen[84]/VPB
+ ANTENNA_mprj_la_oen[84]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[67] la_oen[67] ANTENNA_mprj_la_oen[67]/VGND VSUBS ANTENNA_mprj_la_oen[67]/VPB
+ ANTENNA_mprj_la_oen[67]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[4] wbs_dat_i[4] ANTENNA_mprj_wbs_dat_i[4]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[4]/VPB
+ ANTENNA_mprj_wbs_dat_i[4]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[3] wbs_adr_i[3] ANTENNA_mprj_wbs_adr_i[3]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[3]/VPB
+ ANTENNA_mprj_wbs_adr_i[3]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[101] la_data_in[101] ANTENNA_mprj_la_data_in[101]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[101]/VPB ANTENNA_mprj_la_data_in[101]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[31] la_data_in[31] ANTENNA_mprj_la_data_in[31]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[31]/VPB ANTENNA_mprj_la_data_in[31]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[14] la_data_in[14] ANTENNA_mprj_la_data_in[14]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[14]/VPB ANTENNA_mprj_la_data_in[14]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[126] la_oen[126] ANTENNA_mprj_la_oen[126]/VGND VSUBS ANTENNA_mprj_la_oen[126]/VPB
+ ANTENNA_mprj_la_oen[126]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[109] la_oen[109] ANTENNA_mprj_la_oen[109]/VGND VSUBS ANTENNA_mprj_la_oen[109]/VPB
+ ANTENNA_mprj_la_oen[109]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[83] la_oen[83] ANTENNA_mprj_la_oen[83]/VGND VSUBS ANTENNA_mprj_la_oen[83]/VPB
+ ANTENNA_mprj_la_oen[83]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[11] wbs_adr_i[11] ANTENNA_mprj_wbs_adr_i[11]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[11]/VPB
+ ANTENNA_mprj_wbs_adr_i[11]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[24] wbs_dat_i[24] ANTENNA_mprj_wbs_dat_i[24]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[24]/VPB
+ ANTENNA_mprj_wbs_dat_i[24]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[6] la_oen[6] ANTENNA_mprj_la_oen[6]/VGND VSUBS ANTENNA_mprj_la_oen[6]/VPB
+ ANTENNA_mprj_la_oen[6]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[66] la_oen[66] ANTENNA_mprj_la_oen[66]/VGND VSUBS ANTENNA_mprj_la_oen[66]/VPB
+ ANTENNA_mprj_la_oen[66]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_adr_i[2] wbs_adr_i[2] ANTENNA_mprj_wbs_adr_i[2]/VGND VSUBS ANTENNA_mprj_wbs_adr_i[2]/VPB
+ ANTENNA_mprj_wbs_adr_i[2]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_dat_i[3] wbs_dat_i[3] ANTENNA_mprj_wbs_dat_i[3]/VGND VSUBS ANTENNA_mprj_wbs_dat_i[3]/VPB
+ ANTENNA_mprj_wbs_dat_i[3]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_wbs_sel_i[3] wbs_sel_i[3] ANTENNA_mprj_wbs_sel_i[3]/VGND VSUBS ANTENNA_mprj_wbs_sel_i[3]/VPB
+ ANTENNA_mprj_wbs_sel_i[3]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_oen[49] la_oen[49] ANTENNA_mprj_la_oen[49]/VGND VSUBS ANTENNA_mprj_la_oen[49]/VPB
+ ANTENNA_mprj_la_oen[49]/VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_la_data_in[30] la_data_in[30] ANTENNA_mprj_la_data_in[30]/VGND VSUBS
+ ANTENNA_mprj_la_data_in[30]/VPB ANTENNA_mprj_la_data_in[30]/VPWR sky130_fd_sc_hd__diode_2
.ends

